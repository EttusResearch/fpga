//////////////////////////////////////
//
//  2017 Ettus Research
//
//////////////////////////////////////

module n310_tx_frontend
(

  input [31:0] tx_in,
  output [31:0] tx_out
);

assign tx_out = tx_in;

endmodule
