//////////////////////////////////////
//
//  2017 Ettus Research
//
//////////////////////////////////////

module n310_rx_frontend
(

  input [31:0] rx_in,
  output [31:0] rx_out
);

assign rx_out = rx_in;

endmodule
