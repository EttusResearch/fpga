/////////////////////////////////////////////////////////////////////
//
// Copyright 2016-2017 Ettus Research
//
// N3xx TOP
//
// Rev C Brimstone MB
//
// Rev C Magnesium DB
//
//////////////////////////////////////////////////////////////////////

module n310
(

   inout [11:0] FPGA_GPIO,

   input FPGA_REFCLK_P,
   input FPGA_REFCLK_N,
   input REF_1PPS_IN,
   //input REF_1PPS_IN_MGMT,
   output REF_1PPS_OUT,

   //TDC
   inout aUnusedPinForTdcA0,
   inout aUnusedPinForTdcA1,
   inout aUnusedPinForTdcB0,
   inout aUnusedPinForTdcB1,

   //input NPIO_0_RX0_P,
   //input NPIO_0_RX0_N,
   //input NPIO_0_RX1_P,
   //input NPIO_0_RX1_N,
   //output NPIO_0_TX0_P,
   //output NPIO_0_TX0_N,
   //output NPIO_0_TX1_P,
   //output NPIO_0_TX1_N,
   //input NPIO_1_RX0_P,
   //input NPIO_1_RX0_N,
   //input NPIO_1_RX1_P,
   //input NPIO_1_RX1_N,
   //output NPIO_1_TX0_P,
   //output NPIO_1_TX0_N,
   //output NPIO_1_TX1_P,
   //output NPIO_1_TX1_N,
   //input NPIO_2_RX0_P,
   //input NPIO_2_RX0_N,
   //input NPIO_2_RX1_P,
   //input NPIO_2_RX1_N,
   //output NPIO_2_TX0_P,
   //output NPIO_2_TX0_N,
   //output NPIO_2_TX1_P,
   //output NPIO_2_TX1_N,
   //TODO: Uncomment when connected here
   //input NPIO_0_RXSYNC_0_P, NPIO_0_RXSYNC_1_P,
   //input NPIO_0_RXSYNC_0_N, NPIO_0_RXSYNC_1_N,
   //output NPIO_0_TXSYNC_0_P, NPIO_0_TXSYNC_1_P,
   //output NPIO_0_TXSYNC_0_N, NPIO_0_TXSYNC_1_N,
   //input NPIO_1_RXSYNC_0_P, NPIO_1_RXSYNC_1_P,
   //input NPIO_1_RXSYNC_0_N, NPIO_1_RXSYNC_1_N,
   //output NPIO_1_TXSYNC_0_P, NPIO_1_TXSYNC_1_P,
   //output NPIO_1_TXSYNC_0_N, NPIO_1_TXSYNC_1_N,
   //input NPIO_2_RXSYNC_0_P, NPIO_2_RXSYNC_1_P,
   //input NPIO_2_RXSYNC_0_N, NPIO_2_RXSYNC_1_N,
   //output NPIO_2_TXSYNC_0_P, NPIO_2_TXSYNC_1_P,
   //output NPIO_2_TXSYNC_0_N, NPIO_2_TXSYNC_1_N,

   //GPS
   input GPS_1PPS,
   //input GPS_1PPS_RAW,

   //Misc
   input ENET0_CLK125,
   //inout ENET0_PTP,
   //output ENET0_PTP_DIR,
   //inout ATSHA204_SDA,
   input FPGA_PL_RESETN, // TODO:  Add to reset logic
   output reg [1:0] FPGA_TEST,
   //input PWR_CLK_FPGA, // TODO: check direction

   //White Rabbit
   //input WB_20MHZ_P,
   //input WB_20MHZ_N,
   //output WB_DAC_DIN,
   //output WB_DAC_NCLR,
   //output WB_DAC_NLDAC,
   //output WB_DAC_NSYNC,
   //output WB_DAC_SCLK,
   //output PWREN_CLK_WB_20MHZ,

   //LEDS
   output PANEL_LED_GPS,
   output PANEL_LED_LINK,
   output PANEL_LED_PPS,
   output PANEL_LED_REF,

   // ARM Connections
   inout [53:0]  MIO,
   input         PS_SRSTB,
   input         PS_CLK,
   input         PS_PORB,
   inout         DDR_Clk,
   inout         DDR_Clk_n,
   inout         DDR_CKE,
   inout         DDR_CS_n,
   inout         DDR_RAS_n,
   inout         DDR_CAS_n,
   inout         DDR_WEB,
   inout [2:0]   DDR_BankAddr,
   inout [14:0]  DDR_Addr,
   inout         DDR_ODT,
   inout         DDR_DRSTB,
   inout [31:0]  DDR_DQ,
   inout [3:0]   DDR_DM,
   inout [3:0]   DDR_DQS,
   inout [3:0]   DDR_DQS_n,
   inout         DDR_VRP,
   inout         DDR_VRN,


   ///////////////////////////////////
   //
   // High Speed SPF+ signals and clocking
   //
   ///////////////////////////////////

   //input WB_CDCM_CLK1_P,
   //input WB_CDCM_CLK1_N,

`ifdef BUILD_1G
   input WB_CDCM_CLK2_P,
   input WB_CDCM_CLK2_N,
`endif

`ifdef BUILD_10G
   input MGT156MHZ_CLK1_P,
   input MGT156MHZ_CLK1_N,
`endif
`ifdef BUILD_AURORA
   input MGT156MHZ_CLK1_P,
   input MGT156MHZ_CLK1_N,
`endif

   input SFP_0_RX_P, input SFP_0_RX_N,
   output SFP_0_TX_P, output SFP_0_TX_N,
   input SFP_1_RX_P, input SFP_1_RX_N,
   output SFP_1_TX_P, output SFP_1_TX_N,


   ///////////////////////////////////
   //
   // DRAM Interface
   //
   ///////////////////////////////////
   inout [31:0] ddr3_dq,     // Data pins. Input for Reads, Output for Writes.
   inout [3:0] ddr3_dqs_n,   // Data Strobes. Input for Reads, Output for Writes.
   inout [3:0] ddr3_dqs_p,
   //
   output [15:0] ddr3_addr,  // Address
   output [2:0] ddr3_ba,     // Bank Address
   output ddr3_ras_n,        // Row Address Strobe.
   output ddr3_cas_n,        // Column address select
   output ddr3_we_n,         // Write Enable
   output ddr3_reset_n,      // SDRAM reset pin.
   output [0:0] ddr3_ck_p,         // Differential clock
   output [0:0] ddr3_ck_n,
   output [0:0] ddr3_cke,    // Clock Enable
   output [0:0] ddr3_cs_n,         // Chip Select
   output [3:0] ddr3_dm,     // Data Mask [3] = UDM.U26, [2] = LDM.U26, ...
   output [0:0] ddr3_odt,    // On-Die termination enable.
   //
   input sys_clk_p,          // Differential
   input sys_clk_n,          // 100MHz clock source to generate DDR3 clocking.


   ///////////////////////////////////
   //
   // Supporting I/O for SPF+ interfaces
   //  (non high speed stuff)
   //
   ///////////////////////////////////

   //SFP+ 0, Slow Speed, Bank 13 3.3V
   //input SFP_0_I2C_NPRESENT,
   output SFP_0_LED_A,
   output SFP_0_LED_B,
   input SFP_0_LOS,
   output SFP_0_RS0,
   output SFP_0_RS1,
   output SFP_0_TXDISABLE,
   input SFP_0_TXFAULT,

   //SFP+ 1, Slow Speed, Bank 13 3.3V
   //input SFP_1_I2C_NPRESENT,
   output SFP_1_LED_A,
   output SFP_1_LED_B,
   input SFP_1_LOS,
   output SFP_1_RS0,
   output SFP_1_RS1,
   output SFP_1_TXDISABLE,
   input SFP_1_TXFAULT,

   //USRP IO A
   output        DBA_CPLD_PS_SPI_SCLK,
   output        DBA_CPLD_PS_SPI_LE,
   output        DBA_CPLD_PS_SPI_SDI,
   input         DBA_CPLD_PS_SPI_SDO,
   output [1:0]  DBA_CPLD_PS_SPI_ADDR,

   output        DBA_ATR_RX_1,
   output        DBA_ATR_RX_2,
   output        DBA_ATR_TX_1,
   output        DBA_ATR_TX_2,

   output [5:0]  DBA_CH1_TX_DSA_DATA,
   output [5:0]  DBA_CH1_RX_DSA_DATA,
   output [5:0]  DBA_CH2_TX_DSA_DATA,
   output [5:0]  DBA_CH2_RX_DSA_DATA,

   output        DBA_CPLD_PL_SPI_SCLK,
   output        DBA_CPLD_PL_SPI_LE,
   output        DBA_CPLD_PL_SPI_SDI,
   input         DBA_CPLD_PL_SPI_SDO,
   output [2:0]  DBA_CPLD_PL_SPI_ADDR,

   output        DBA_MYK_SPI_SCLK,
   output        DBA_MYK_SPI_CS_n,
   input         DBA_MYK_SPI_SDO,
   output        DBA_MYK_SPI_SDIO,
   input         DBA_MYK_INTRQ,

   output        DBA_MYK_SYNC_IN_n,
   input         DBA_MYK_SYNC_OUT_n,

   output        DBA_CPLD_JTAG_TCK,
   output        DBA_CPLD_JTAG_TMS,
   output        DBA_CPLD_JTAG_TDI,
   input         DBA_CPLD_JTAG_TDO,

   output        DBA_MYK_GPIO_0,
   output        DBA_MYK_GPIO_1,
   output        DBA_MYK_GPIO_3,
   output        DBA_MYK_GPIO_4,
   output        DBA_MYK_GPIO_12,
   output        DBA_MYK_GPIO_13,
   output        DBA_MYK_GPIO_14,
   output        DBA_MYK_GPIO_15,

   input         DBA_FPGA_CLK_p,
   input         DBA_FPGA_CLK_n,
   input         DBA_FPGA_SYSREF_p,
   input         DBA_FPGA_SYSREF_n,

   input         USRPIO_A_MGTCLK_P,
   input         USRPIO_A_MGTCLK_N,

   input  [3:0]  USRPIO_A_RX_P,
   input  [3:0]  USRPIO_A_RX_N,
   output [3:0]  USRPIO_A_TX_P,
   output [3:0]  USRPIO_A_TX_N,


   //USRP IO B
   output        DBB_CPLD_PS_SPI_SCLK,
   output        DBB_CPLD_PS_SPI_LE,
   output        DBB_CPLD_PS_SPI_SDI,
   input         DBB_CPLD_PS_SPI_SDO,
   output [1:0]  DBB_CPLD_PS_SPI_ADDR,

   output        DBB_ATR_RX_1,
   output        DBB_ATR_RX_2,
   output        DBB_ATR_TX_1,
   output        DBB_ATR_TX_2,

   output [5:0]  DBB_CH1_TX_DSA_DATA,
   output [5:0]  DBB_CH1_RX_DSA_DATA,
   output [5:0]  DBB_CH2_TX_DSA_DATA,
   output [5:0]  DBB_CH2_RX_DSA_DATA,

   output        DBB_CPLD_PL_SPI_SCLK,
   output        DBB_CPLD_PL_SPI_LE,
   output        DBB_CPLD_PL_SPI_SDI,
   input         DBB_CPLD_PL_SPI_SDO,
   output [2:0]  DBB_CPLD_PL_SPI_ADDR,

   output        DBB_MYK_SPI_SCLK,
   output        DBB_MYK_SPI_CS_n,
   input         DBB_MYK_SPI_SDO,
   output        DBB_MYK_SPI_SDIO,
   input         DBB_MYK_INTRQ,

   output        DBB_MYK_SYNC_IN_n,
   input         DBB_MYK_SYNC_OUT_n,

   output        DBB_CPLD_JTAG_TCK,
   output        DBB_CPLD_JTAG_TMS,
   output        DBB_CPLD_JTAG_TDI,
   input         DBB_CPLD_JTAG_TDO,

   output        DBB_MYK_GPIO_0,
   output        DBB_MYK_GPIO_1,
   output        DBB_MYK_GPIO_3,
   output        DBB_MYK_GPIO_4,
   output        DBB_MYK_GPIO_12,
   output        DBB_MYK_GPIO_13,
   output        DBB_MYK_GPIO_14,
   output        DBB_MYK_GPIO_15,

   input         DBB_FPGA_CLK_p,
   input         DBB_FPGA_CLK_n,
   input         DBB_FPGA_SYSREF_p,
   input         DBB_FPGA_SYSREF_n,

   input         USRPIO_B_MGTCLK_P,
   input         USRPIO_B_MGTCLK_N,

   input  [3:0]  USRPIO_B_RX_P,
   input  [3:0]  USRPIO_B_RX_N,
   output [3:0]  USRPIO_B_TX_P,
   output [3:0]  USRPIO_B_TX_N




);

  localparam N_AXILITE_SLAVES = 4;
  localparam REG_AWIDTH = 14; // log2(0x4000)
  localparam REG_DWIDTH = 32;

  // TODO: Add sw_rst
  wire bus_clk;
  wire bus_rst;
  wire global_rst;

  // Internal connections to PS
  // HP0 -- High Performance port 0, FPGA is the master
  wire [5:0]  S_AXI_HP0_AWID;
  wire [31:0] S_AXI_HP0_AWADDR;
  wire [2:0]  S_AXI_HP0_AWPROT;
  wire        S_AXI_HP0_AWVALID;
  wire        S_AXI_HP0_AWREADY;
  wire [63:0] S_AXI_HP0_WDATA;
  wire [7:0]  S_AXI_HP0_WSTRB;
  wire        S_AXI_HP0_WVALID;
  wire        S_AXI_HP0_WREADY;
  wire [1:0]  S_AXI_HP0_BRESP;
  wire        S_AXI_HP0_BVALID;
  wire        S_AXI_HP0_BREADY;
  wire [5:0]  S_AXI_HP0_ARID;
  wire [31:0] S_AXI_HP0_ARADDR;
  wire [2:0]  S_AXI_HP0_ARPROT;
  wire        S_AXI_HP0_ARVALID;
  wire        S_AXI_HP0_ARREADY;
  wire [63:0] S_AXI_HP0_RDATA;
  wire [1:0]  S_AXI_HP0_RRESP;
  wire        S_AXI_HP0_RVALID;
  wire        S_AXI_HP0_RREADY;
  wire [3:0]  S_AXI_HP0_ARCACHE;
  wire [7:0]  S_AXI_HP0_AWLEN;
  wire [2:0]  S_AXI_HP0_AWSIZE;
  wire [1:0]  S_AXI_HP0_AWBURST;
  wire [3:0]  S_AXI_HP0_AWCACHE;
  wire        S_AXI_HP0_WLAST;
  wire [7:0]  S_AXI_HP0_ARLEN;
  wire [1:0]  S_AXI_HP0_ARBURST;
  wire [2:0]  S_AXI_HP0_ARSIZE;

  // GP0 -- General Purpose port 0, FPGA is the master
  wire [5:0]  S_AXI_GP0_AWID;
  wire [31:0] S_AXI_GP0_AWADDR;
  wire [2:0]  S_AXI_GP0_AWPROT;
  wire        S_AXI_GP0_AWVALID;
  wire        S_AXI_GP0_AWREADY;
  wire [31:0] S_AXI_GP0_WDATA;
  wire [3:0]  S_AXI_GP0_WSTRB;
  wire        S_AXI_GP0_WVALID;
  wire        S_AXI_GP0_WREADY;
  wire [1:0]  S_AXI_GP0_BRESP;
  wire        S_AXI_GP0_BVALID;
  wire        S_AXI_GP0_BREADY;
  wire [5:0]  S_AXI_GP0_ARID;
  wire [31:0] S_AXI_GP0_ARADDR;
  wire [2:0]  S_AXI_GP0_ARPROT;
  wire        S_AXI_GP0_ARVALID;
  wire        S_AXI_GP0_ARREADY;
  wire [31:0] S_AXI_GP0_RDATA;
  wire [1:0]  S_AXI_GP0_RRESP;
  wire        S_AXI_GP0_RVALID;
  wire        S_AXI_GP0_RREADY;
  wire [3:0]  S_AXI_GP0_ARCACHE;
  wire [7:0]  S_AXI_GP0_AWLEN;
  wire [2:0]  S_AXI_GP0_AWSIZE;
  wire [1:0]  S_AXI_GP0_AWBURST;
  wire [3:0]  S_AXI_GP0_AWCACHE;
  wire        S_AXI_GP0_WLAST;
  wire [7:0]  S_AXI_GP0_ARLEN;
  wire [1:0]  S_AXI_GP0_ARBURST;
  wire [2:0]  S_AXI_GP0_ARSIZE;

  // HP1 -- High Performance port 1, FPGA is the master
  wire [5:0]  S_AXI_HP1_AWID;
  wire [31:0] S_AXI_HP1_AWADDR;
  wire [2:0]  S_AXI_HP1_AWPROT;
  wire        S_AXI_HP1_AWVALID;
  wire        S_AXI_HP1_AWREADY;
  wire [63:0] S_AXI_HP1_WDATA;
  wire [7:0]  S_AXI_HP1_WSTRB;
  wire        S_AXI_HP1_WVALID;
  wire        S_AXI_HP1_WREADY;
  wire [1:0]  S_AXI_HP1_BRESP;
  wire        S_AXI_HP1_BVALID;
  wire        S_AXI_HP1_BREADY;
  wire [5:0]  S_AXI_HP1_ARID;
  wire [31:0] S_AXI_HP1_ARADDR;
  wire [2:0]  S_AXI_HP1_ARPROT;
  wire        S_AXI_HP1_ARVALID;
  wire        S_AXI_HP1_ARREADY;
  wire [63:0] S_AXI_HP1_RDATA;
  wire [1:0]  S_AXI_HP1_RRESP;
  wire        S_AXI_HP1_RVALID;
  wire        S_AXI_HP1_RREADY;
  wire [3:0]  S_AXI_HP1_ARCACHE;
  wire [7:0]  S_AXI_HP1_AWLEN;
  wire [2:0]  S_AXI_HP1_AWSIZE;
  wire [1:0]  S_AXI_HP1_AWBURST;
  wire [3:0]  S_AXI_HP1_AWCACHE;
  wire        S_AXI_HP1_WLAST;
  wire [7:0]  S_AXI_HP1_ARLEN;
  wire [1:0]  S_AXI_HP1_ARBURST;
  wire [2:0]  S_AXI_HP1_ARSIZE;

  // GP1 -- General Purpose port 1, FPGA is the master
  wire [5:0]  S_AXI_GP1_AWID;
  wire [31:0] S_AXI_GP1_AWADDR;
  wire [2:0]  S_AXI_GP1_AWPROT;
  wire        S_AXI_GP1_AWVALID;
  wire        S_AXI_GP1_AWREADY;
  wire [31:0] S_AXI_GP1_WDATA;
  wire [3:0]  S_AXI_GP1_WSTRB;
  wire        S_AXI_GP1_WVALID;
  wire        S_AXI_GP1_WREADY;
  wire [1:0]  S_AXI_GP1_BRESP;
  wire        S_AXI_GP1_BVALID;
  wire        S_AXI_GP1_BREADY;
  wire [5:0]  S_AXI_GP1_ARID;
  wire [31:0] S_AXI_GP1_ARADDR;
  wire [2:0]  S_AXI_GP1_ARPROT;
  wire        S_AXI_GP1_ARVALID;
  wire        S_AXI_GP1_ARREADY;
  wire [31:0] S_AXI_GP1_RDATA;
  wire [1:0]  S_AXI_GP1_RRESP;
  wire        S_AXI_GP1_RVALID;
  wire        S_AXI_GP1_RREADY;
  wire [3:0]  S_AXI_GP1_ARCACHE;
  wire [7:0]  S_AXI_GP1_AWLEN;
  wire [2:0]  S_AXI_GP1_AWSIZE;
  wire [1:0]  S_AXI_GP1_AWBURST;
  wire [3:0]  S_AXI_GP1_AWCACHE;
  wire        S_AXI_GP1_WLAST;
  wire [7:0]  S_AXI_GP1_ARLEN;
  wire [1:0]  S_AXI_GP1_ARBURST;
  wire [2:0]  S_AXI_GP1_ARSIZE;

  // GP0 -- General Purpose port 0, FPGA is the slave
  wire        M_AXI_GP0_ARVALID;
  wire        M_AXI_GP0_AWVALID;
  wire        M_AXI_GP0_BREADY;
  wire        M_AXI_GP0_RREADY;
  wire        M_AXI_GP0_WVALID;
  wire [11:0] M_AXI_GP0_ARID;
  wire [11:0] M_AXI_GP0_AWID;
  wire [11:0] M_AXI_GP0_WID;
  wire [31:0] M_AXI_GP0_ARADDR;
  wire [31:0] M_AXI_GP0_AWADDR;
  wire [31:0] M_AXI_GP0_WDATA;
  wire [3:0]  M_AXI_GP0_WSTRB;
  wire        M_AXI_GP0_ARREADY;
  wire        M_AXI_GP0_AWREADY;
  wire        M_AXI_GP0_BVALID;
  wire        M_AXI_GP0_RLAST;
  wire        M_AXI_GP0_RVALID;
  wire        M_AXI_GP0_WREADY;
  wire [1:0]  M_AXI_GP0_BRESP;
  wire [1:0]  M_AXI_GP0_RRESP;
  wire [31:0] M_AXI_GP0_RDATA;

  wire        M_AXI_GP0_ARVALID_S0;
  wire        M_AXI_GP0_AWVALID_S0;
  wire        M_AXI_GP0_BREADY_S0;
  wire        M_AXI_GP0_RREADY_S0;
  wire        M_AXI_GP0_WVALID_S0;
  wire [11:0] M_AXI_GP0_ARID_S0;
  wire [11:0] M_AXI_GP0_AWID_S0;
  wire [11:0] M_AXI_GP0_WID_S0;
  wire [31:0] M_AXI_GP0_ARADDR_S0;
  wire [31:0] M_AXI_GP0_AWADDR_S0;
  wire [31:0] M_AXI_GP0_WDATA_S0;
  wire [3:0]  M_AXI_GP0_WSTRB_S0;
  wire        M_AXI_GP0_ARREADY_S0;
  wire        M_AXI_GP0_AWREADY_S0;
  wire        M_AXI_GP0_BVALID_S0;
  wire        M_AXI_GP0_RLAST_S0;
  wire        M_AXI_GP0_RVALID_S0;
  wire        M_AXI_GP0_WREADY_S0;
  wire [1:0]  M_AXI_GP0_BRESP_S0;
  wire [1:0]  M_AXI_GP0_RRESP_S0;
  wire [31:0] M_AXI_GP0_RDATA_S0;

  wire        M_AXI_GP0_ARVALID_S1;
  wire        M_AXI_GP0_AWVALID_S1;
  wire        M_AXI_GP0_BREADY_S1;
  wire        M_AXI_GP0_RREADY_S1;
  wire        M_AXI_GP0_WVALID_S1;
  wire [11:0] M_AXI_GP0_ARID_S1;
  wire [11:0] M_AXI_GP0_AWID_S1;
  wire [11:0] M_AXI_GP0_WID_S1;
  wire [31:0] M_AXI_GP0_ARADDR_S1;
  wire [31:0] M_AXI_GP0_AWADDR_S1;
  wire [31:0] M_AXI_GP0_WDATA_S1;
  wire [3:0]  M_AXI_GP0_WSTRB_S1;
  wire        M_AXI_GP0_ARREADY_S1;
  wire        M_AXI_GP0_AWREADY_S1;
  wire        M_AXI_GP0_BVALID_S1;
  wire        M_AXI_GP0_RLAST_S1;
  wire        M_AXI_GP0_RVALID_S1;
  wire        M_AXI_GP0_WREADY_S1;
  wire [1:0]  M_AXI_GP0_BRESP_S1;
  wire [1:0]  M_AXI_GP0_RRESP_S1;
  wire [31:0] M_AXI_GP0_RDATA_S1;

  wire        M_AXI_GP0_ARVALID_S2;
  wire        M_AXI_GP0_AWVALID_S2;
  wire        M_AXI_GP0_BREADY_S2;
  wire        M_AXI_GP0_RREADY_S2;
  wire        M_AXI_GP0_WVALID_S2;
  wire [11:0] M_AXI_GP0_ARID_S2;
  wire [11:0] M_AXI_GP0_AWID_S2;
  wire [11:0] M_AXI_GP0_WID_S2;
  wire [31:0] M_AXI_GP0_ARADDR_S2;
  wire [31:0] M_AXI_GP0_AWADDR_S2;
  wire [31:0] M_AXI_GP0_WDATA_S2;
  wire [3:0]  M_AXI_GP0_WSTRB_S2;
  wire        M_AXI_GP0_ARREADY_S2;
  wire        M_AXI_GP0_AWREADY_S2;
  wire        M_AXI_GP0_BVALID_S2;
  wire        M_AXI_GP0_RLAST_S2;
  wire        M_AXI_GP0_RVALID_S2;
  wire        M_AXI_GP0_WREADY_S2;
  wire [1:0]  M_AXI_GP0_BRESP_S2;
  wire [1:0]  M_AXI_GP0_RRESP_S2;
  wire [31:0] M_AXI_GP0_RDATA_S2;

  wire        M_AXI_GP0_ARVALID_S3;
  wire        M_AXI_GP0_AWVALID_S3;
  wire        M_AXI_GP0_BREADY_S3;
  wire        M_AXI_GP0_RREADY_S3;
  wire        M_AXI_GP0_WVALID_S3;
  wire [11:0] M_AXI_GP0_ARID_S3;
  wire [11:0] M_AXI_GP0_AWID_S3;
  wire [11:0] M_AXI_GP0_WID_S3;
  wire [31:0] M_AXI_GP0_ARADDR_S3;
  wire [31:0] M_AXI_GP0_AWADDR_S3;
  wire [31:0] M_AXI_GP0_WDATA_S3;
  wire [3:0]  M_AXI_GP0_WSTRB_S3;
  wire        M_AXI_GP0_ARREADY_S3;
  wire        M_AXI_GP0_AWREADY_S3;
  wire        M_AXI_GP0_BVALID_S3;
  wire        M_AXI_GP0_RLAST_S3;
  wire        M_AXI_GP0_RVALID_S3;
  wire        M_AXI_GP0_WREADY_S3;
  wire [1:0]  M_AXI_GP0_BRESP_S3;
  wire [1:0]  M_AXI_GP0_RRESP_S3;
  wire [31:0] M_AXI_GP0_RDATA_S3;

  wire        M_AXI_GP0_ARVALID_S4;
  wire        M_AXI_GP0_AWVALID_S4;
  wire        M_AXI_GP0_BREADY_S4;
  wire        M_AXI_GP0_RREADY_S4;
  wire        M_AXI_GP0_WVALID_S4;
  wire [11:0] M_AXI_GP0_ARID_S4;
  wire [11:0] M_AXI_GP0_AWID_S4;
  wire [11:0] M_AXI_GP0_WID_S4;
  wire [31:0] M_AXI_GP0_ARADDR_S4;
  wire [31:0] M_AXI_GP0_AWADDR_S4;
  wire [31:0] M_AXI_GP0_WDATA_S4;
  wire [3:0]  M_AXI_GP0_WSTRB_S4;
  wire        M_AXI_GP0_ARREADY_S4;
  wire        M_AXI_GP0_AWREADY_S4;
  wire        M_AXI_GP0_BVALID_S4;
  wire        M_AXI_GP0_RLAST_S4;
  wire        M_AXI_GP0_RVALID_S4;
  wire        M_AXI_GP0_WREADY_S4;
  wire [1:0]  M_AXI_GP0_BRESP_S4;
  wire [1:0]  M_AXI_GP0_RRESP_S4;
  wire [31:0] M_AXI_GP0_RDATA_S4;

  wire        M_AXI_GP0_ARVALID_S5;
  wire        M_AXI_GP0_AWVALID_S5;
  wire        M_AXI_GP0_BREADY_S5;
  wire        M_AXI_GP0_RREADY_S5;
  wire        M_AXI_GP0_WVALID_S5;
  wire [11:0] M_AXI_GP0_ARID_S5;
  wire [11:0] M_AXI_GP0_AWID_S5;
  wire [11:0] M_AXI_GP0_WID_S5;
  wire [31:0] M_AXI_GP0_ARADDR_S5;
  wire [31:0] M_AXI_GP0_AWADDR_S5;
  wire [31:0] M_AXI_GP0_WDATA_S5;
  wire [3:0]  M_AXI_GP0_WSTRB_S5;
  wire        M_AXI_GP0_ARREADY_S5;
  wire        M_AXI_GP0_AWREADY_S5;
  wire        M_AXI_GP0_BVALID_S5;
  wire        M_AXI_GP0_RLAST_S5;
  wire        M_AXI_GP0_RVALID_S5;
  wire        M_AXI_GP0_WREADY_S5;
  wire [1:0]  M_AXI_GP0_BRESP_S5;
  wire [1:0]  M_AXI_GP0_RRESP_S5;
  wire [31:0] M_AXI_GP0_RDATA_S5;

  wire        M_AXI_GP0_ARVALID_S6;
  wire        M_AXI_GP0_AWVALID_S6;
  wire        M_AXI_GP0_BREADY_S6;
  wire        M_AXI_GP0_RREADY_S6;
  wire        M_AXI_GP0_WVALID_S6;
  wire [11:0] M_AXI_GP0_ARID_S6;
  wire [11:0] M_AXI_GP0_AWID_S6;
  wire [11:0] M_AXI_GP0_WID_S6;
  wire [31:0] M_AXI_GP0_ARADDR_S6;
  wire [31:0] M_AXI_GP0_AWADDR_S6;
  wire [31:0] M_AXI_GP0_WDATA_S6;
  wire [3:0]  M_AXI_GP0_WSTRB_S6;
  wire        M_AXI_GP0_ARREADY_S6;
  wire        M_AXI_GP0_AWREADY_S6;
  wire        M_AXI_GP0_BVALID_S6;
  wire        M_AXI_GP0_RLAST_S6;
  wire        M_AXI_GP0_RVALID_S6;
  wire        M_AXI_GP0_WREADY_S6;
  wire [1:0]  M_AXI_GP0_BRESP_S6;
  wire [1:0]  M_AXI_GP0_RRESP_S6;
  wire [31:0] M_AXI_GP0_RDATA_S6;

  wire        M_AXI_GP0_ARVALID_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_AWVALID_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_BREADY_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_RREADY_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_WVALID_S[N_AXILITE_SLAVES-1:0];
  wire [11:0] M_AXI_GP0_ARID_S[N_AXILITE_SLAVES-1:0];
  wire [11:0] M_AXI_GP0_AWID_S[N_AXILITE_SLAVES-1:0];
  wire [11:0] M_AXI_GP0_WID_S[N_AXILITE_SLAVES-1:0];
  wire [31:0] M_AXI_GP0_ARADDR_S[N_AXILITE_SLAVES-1:0];
  wire [31:0] M_AXI_GP0_AWADDR_S[N_AXILITE_SLAVES-1:0];
  wire [31:0] M_AXI_GP0_WDATA_S[N_AXILITE_SLAVES-1:0];
  wire [3:0]  M_AXI_GP0_WSTRB_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_ARREADY_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_AWREADY_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_BVALID_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_RLAST_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_RVALID_S[N_AXILITE_SLAVES-1:0];
  wire        M_AXI_GP0_WREADY_S[N_AXILITE_SLAVES-1:0];
  wire [1:0]  M_AXI_GP0_BRESP_S[N_AXILITE_SLAVES-1:0];
  wire [1:0]  M_AXI_GP0_RRESP_S[N_AXILITE_SLAVES-1:0];
  wire [31:0] M_AXI_GP0_RDATA_S[N_AXILITE_SLAVES-1:0];

  wire [15:0] IRQ_F2P;
  wire        clk100;
  wire        clk40;
  wire        FCLK_RESET0;
  wire        FCLK_RESET0N = ~FCLK_RESET0;

  wire [1:0] USB0_PORT_INDCTL;
  wire       USB0_VBUS_PWRSELECT;
  wire       USB0_VBUS_PWRFAULT;

  /////////////////////////////////////////////////////////////////////
  //
  // power-on-reset logic.
  //
  //////////////////////////////////////////////////////////////////////
  por_gen por_gen(.clk(bus_clk), .reset_out(global_rst));

  //////////////////////////////////////////////////////////////////////
  //
  // Configure SFP+ clocking
  //
  //////////////////////////////////////////////////////////////////////
  //
  //   PL Clocks : ---------------------------------------------------------------------------
  //   xgige_refclk (156): MGT156MHZ_CLK1_P > GTX IBUF > IBUFDS_GTE2  > xgige_refclk
  //   clk156            : MGT156MHZ_CLK1_P > GTX IBUF > IBUFDS_GTE2  > BUFG  > clk156
  //   gige_refclk (125) : WB_CDCM_CLK2_P   > GTX IBUF > IBUFDS_GTE2  > gige_refclk
  //   gige_refclk_bufg  : WB_CDCM_CLK2_P   > GTX IBUF > IBUFDS_GTE2  > gige_refclk_bufg
  //   RefClk (10)       : FPGA_REFCLK_P    >   IBUFDS > ref_clk
  //
  //   PS Clocks to PL:
  //   FCLK_CLK0 :      100 MHz
  //   FCLK_CLK1 :       40 MHz
  //   FCLK_CLK2 : 166.6667 MHz
  //   FCLK_CLK3 :      200 MHz
  //
  /////////////////////////////////////////////////////////////////////

  /////////////////////////////////////////////////////////////////////
  //
  // 10MHz Reference clock
  //
  //////////////////////////////////////////////////////////////////////

  wire ref_clk_buf;
  wire ref_clk;

  wire radio_clk;
  wire radio_clkB;
  wire radio_clk_2x;
  wire radio_clk_2xB;

  wire meas_clk_ref;
  wire meas_clk;
  wire meas_clk_reset;
  wire meas_clk_locked;

  // FPGA Reference Clock Buffering
  //
  // Only require an IBUF and BUFG here, since an MMCM is (thankfully) not needed
  // to meet timing with the PPS signal.
  IBUFDS IBUFDS_ref_clk (
       .O(ref_clk_buf),
       .I(FPGA_REFCLK_P),
       .IB(FPGA_REFCLK_N)
   );

  BUFG BUFG_ref_clk (
       .O(ref_clk),
       .I(ref_clk_buf)
   );

  // Measurement Clock MMCM Instantiation
  //
  // This must be an MMCM to hit the weird rates we need for meas_clk.
  MeasClkMmcm MeasClkMmcmx (
    .clk_in1 (meas_clk_ref),
    .clk_out1(meas_clk),
    .reset   (meas_clk_reset),
    .locked  (meas_clk_locked)
  );



  wire radio_rst;

  //FIXME RESET SYNC may need more or'd inputs.
  reset_sync radio_reset_sync (
     .clk(radio_clk),
     .reset_in(global_rst),
     //FIXME EXAMPLE of various reset_in sources
     //.reset_in(global_rst || !bus_clk_locked || sw_rst[1]),
     .reset_out(radio_rst)
  );

  reset_sync int_reset_sync (
     .clk(bus_clk),
     .reset_in(global_rst),
     .reset_out(bus_rst)
  );

`ifdef BUILD_1G
   wire  gige_refclk, gige_refclk_bufg;

   one_gige_phy_clk_gen gige_clk_gen_i (
      .areset(global_rst),
      .refclk_p(WB_CDCM_CLK2_P),
      .refclk_n(WB_CDCM_CLK2_N),
      .refclk(gige_refclk),
      .refclk_bufg(gige_refclk_bufg)
   );

   // FIXME
   assign SFP_0_RS0  = 1'b0;
   assign SFP_0_RS1  = 1'b0;
   assign SFP_1_RS0  = 1'b0;
   assign SFP_1_RS1  = 1'b0;

`endif

`ifdef BUILD_10G
   wire  xgige_refclk;
   wire  xgige_clk156;
   wire  xgige_dclk;

   ten_gige_phy_clk_gen xgige_clk_gen_i (
      .areset(global_rst),
      .refclk_p(MGT156MHZ_CLK1_P),
      .refclk_n(MGT156MHZ_CLK1_N),
      .refclk(xgige_refclk),
      .clk156(xgige_clk156),
      .dclk(xgige_dclk)
   );
   // FIXME
   assign SFP_0_RS0  = 1'b1;
   assign SFP_0_RS1  = 1'b1;
   assign SFP_1_RS0  = 1'b1;
   assign SFP_1_RS1  = 1'b1;

`endif

`ifdef BUILD_AURORA
  wire aurora_refclk, aurora_clk156, aurora_init_clk;
  aurora_phy_clk_gen aurora_clk_gen_i (
    .areset(global_rst),
    .refclk_p(MGT156MHZ_CLK1_P),
    .refclk_n(MGT156MHZ_CLK1_N),
    .refclk(aurora_refclk),
    .clk156(aurora_clk156),
    .init_clk(aurora_init_clk)
  );

   assign SFP_0_RS0  = 1'b1;
   assign SFP_0_RS1  = 1'b1;
   assign SFP_1_RS0  = 1'b1;
   assign SFP_1_RS1  = 1'b1;
`endif

  //If bus_clk freq ever changes, update this paramter accordingly.
  localparam BUS_CLK_RATE = 32'd200000000; //200 MHz bus_clk rate. 

   wire  sfp0_gt_refclk, sfp1_gt_refclk;
   wire  sfp0_gb_refclk, sfp1_gb_refclk;
   wire  sfp0_misc_clk, sfp1_misc_clk;

`ifdef SFP0_10GBE
   assign sfp0_gt_refclk = xgige_refclk;
   assign sfp0_gb_refclk = xgige_clk156;
   assign sfp0_misc_clk  = xgige_dclk;
`endif
`ifdef SFP0_1GBE
   assign sfp0_gt_refclk = gige_refclk;
   assign sfp0_gb_refclk = gige_refclk_bufg;
   assign sfp0_misc_clk  = gige_refclk_bufg;
`endif
`ifdef SFP0_AURORA
   assign sfp0_gt_refclk = aurora_refclk;
   assign sfp0_gb_refclk = aurora_clk156;
   assign sfp0_misc_clk  = aurora_init_clk;
`endif
`ifdef SFP1_10GBE
   assign sfp1_gt_refclk = xgige_refclk;
   assign sfp1_gb_refclk = xgige_clk156;
   assign sfp1_misc_clk  = xgige_dclk;
`endif
`ifdef SFP1_1GBE
   assign sfp1_gt_refclk = gige_refclk;
   assign sfp1_gb_refclk = gige_refclk_bufg;
   assign sfp1_misc_clk  = gige_refclk_bufg;
`endif
`ifdef SFP0_AURORA
   assign sfp1_gt_refclk = aurora_refclk;
   assign sfp1_gb_refclk = aurora_clk156;
   assign sfp1_misc_clk  = aurora_init_clk;
`endif

   wire          gt0_qplloutclk,gt0_qplloutrefclk;
   wire          pma_reset;
   wire          qpllreset;
   wire          qplllock;
   wire          qplloutclk;
   wire          qplloutrefclk;
   wire  [15:0]  sfp0_phy_status;
   wire  [15:0]  sfp1_phy_status;
   wire  [63:0]  e01_tdata, e10_tdata;
   wire  [3:0]   e01_tuser, e10_tuser;
   wire          e01_tlast, e01_tvalid, e01_tready;
   wire          e10_tlast, e10_tvalid, e10_tready;

`ifdef SFP0_1GBE
   //GT COMMON
   one_gig_eth_pcs_pma_gt_common core_gt_common_i
   (
    .GTREFCLK0_IN                (gige_refclk) ,
    .QPLLLOCK_OUT                (),
    .QPLLLOCKDETCLK_IN           (bus_clk),
    .QPLLOUTCLK_OUT              (gt0_qplloutclk),
    .QPLLOUTREFCLK_OUT           (gt0_qplloutrefclk),
    .QPLLREFCLKLOST_OUT          (),
    .QPLLRESET_IN                (pma_reset)
   );
`endif

`ifdef SFP0_10GBE

  // Instantiate the 10GBASER/KR GT Common block
  ten_gig_eth_pcs_pma_gt_common # (
      .WRAPPER_SIM_GTRESET_SPEEDUP("TRUE") ) //Does not affect hardware
  ten_gig_eth_pcs_pma_gt_common_block
    (
     .refclk(xgige_refclk),
     .qpllreset(qpllreset),
     .qplllock(qplllock),
     .qplloutclk(qplloutclk),
     .qplloutrefclk(qplloutrefclk),
     .qpllrefclksel(3'b101 /*GTSOUTHREFCLK0*/)
    );
`endif

`ifdef SFP0_AURORA
  wire qpllrefclklost;

  wire    [7:0]      qpll_drpaddr_in_i = 8'h0;
  wire    [15:0]     qpll_drpdi_in_i = 16'h0;
  wire               qpll_drpen_in_i =  1'b0;
  wire               qpll_drpwe_in_i =  1'b0;
  wire    [15:0]     qpll_drpdo_out_i;
  wire               qpll_drprdy_out_i;

  aurora_64b66b_pcs_pma_gt_common_wrapper gt_common_support (
    .gt_qpllclk_quad1_out      (qplloutclk), //to sfp
    .gt_qpllrefclk_quad1_out   (qplloutrefclk), // to sfp
    .GT0_GTREFCLK0_COMMON_IN   (aurora_refclk),
    //----------------------- Common Block - QPLL Ports ------------------------
    .GT0_QPLLLOCK_OUT          (qplllock), //from 1st sfp
    .GT0_QPLLRESET_IN          (qpllreset), //from 1st sfp
    .GT0_QPLLLOCKDETCLK_IN     (aurora_init_clk),
    .GT0_QPLLREFCLKLOST_OUT    (qpllrefclklost), //from 1st sfp
    //---------------------- Common DRP Ports ---------------------- //not really used???
    .qpll_drpaddr_in           (qpll_drpaddr_in_i),
    .qpll_drpdi_in             (qpll_drpdi_in_i),
    .qpll_drpclk_in            (aurora_init_clk),
    .qpll_drpdo_out            (qpll_drpdo_out_i),
    .qpll_drprdy_out           (qpll_drprdy_out_i),
    .qpll_drpen_in             (qpll_drpen_in_i),
    .qpll_drpwe_in             (qpll_drpwe_in_i)
  );
`endif

  ////////////////////////////////////////////////////////////////////
  // PPS
  // Support for internal or external inputs.
  ///////////////////////////////////////////////////////////////////

  // Generate an internal PPS signal with a 25% duty cycle
  wire r_int_pps;
  pps_generator #(
     .CLK_FREQ(32'd10_000_000), .DUTY_CYCLE(25)
  ) pps_gen (
     .clk(ref_clk), .reset(1'b0), .pps(r_int_pps)
  );

  // PPS MUX - selects internal or external PPS.
  wire [1:0] pps_select;
  wire pps_out_enb;
  reg r_pps_select_ms = 1'b0;
  reg r_pps_select    = 1'b0;
  reg r_pps_ext_ms    = 1'b0;
  reg r_pps_ext       = 1'b0;
  reg pps_refclk      = 1'b0;
  always @(posedge ref_clk) begin

    // Capture the external PPS with a FF before sending to the select. To be safe,
    // we double-synchronize the external signal. If we meet timing (which we should)
    // then this is a two-cycle delay. If we don't meet timing, then it's 1-2 cycles
    // and our system timing is thrown off--but at least our downstream logic doesn't
    // go haywire!
    r_pps_ext_ms <= REF_1PPS_IN;
    r_pps_ext    <= r_pps_ext_ms;

    r_pps_select_ms <= pps_select[0]; // pps_select[1:0] comes from a register in some unknown domain
    r_pps_select    <= r_pps_select_ms;

    if(r_pps_select)
      pps_refclk <= r_int_pps; // pps_select = 1 = internal
    else
      pps_refclk <= r_pps_ext;

    FPGA_TEST[1] <= pps_refclk;
  end

  // PPS out and LED
  assign PANEL_LED_PPS = pps_refclk;


// ARM ethernet 0 bridge signals
  wire [63:0] arm_eth0_tx_tdata;
  wire        arm_eth0_tx_tvalid;
  wire        arm_eth0_tx_tlast;
  wire        arm_eth0_tx_tready;
  wire [3:0]  arm_eth0_tx_tuser;
  wire [7:0]  arm_eth0_tx_tkeep;

  wire [63:0] arm_eth0_tx_tdata_b;
  wire        arm_eth0_tx_tvalid_b;
  wire        arm_eth0_tx_tlast_b;
  wire        arm_eth0_tx_tready_b;
  wire [3:0]  arm_eth0_tx_tuser_b;
  wire [7:0]  arm_eth0_tx_tkeep_b;

  wire [63:0] arm_eth0_rx_tdata;
  wire        arm_eth0_rx_tvalid;
  wire        arm_eth0_rx_tlast;
  wire        arm_eth0_rx_tready;
  wire [3:0]  arm_eth0_rx_tuser;
  wire [7:0]  arm_eth0_rx_tkeep;

  wire [63:0] arm_eth0_rx_tdata_b;
  wire        arm_eth0_rx_tvalid_b;
  wire        arm_eth0_rx_tlast_b;
  wire        arm_eth0_rx_tready_b;
  wire [3:0]  arm_eth0_rx_tuser_b;
  wire [7:0]  arm_eth0_rx_tkeep_b;

  wire        arm_eth0_rx_irq;
  wire        arm_eth0_tx_irq;

  // ARM ethernet 1 bridge signals
  wire [63:0] arm_eth1_tx_tdata;
  wire        arm_eth1_tx_tvalid;
  wire        arm_eth1_tx_tlast;
  wire        arm_eth1_tx_tready;
  wire [3:0]  arm_eth1_tx_tuser;
  wire [7:0]  arm_eth1_tx_tkeep;

  wire [63:0] arm_eth1_tx_tdata_b;
  wire        arm_eth1_tx_tvalid_b;
  wire        arm_eth1_tx_tlast_b;
  wire        arm_eth1_tx_tready_b;
  wire [3:0]  arm_eth1_tx_tuser_b;
  wire [7:0]  arm_eth1_tx_tkeep_b;

  wire [63:0] arm_eth1_rx_tdata;
  wire        arm_eth1_rx_tvalid;
  wire        arm_eth1_rx_tlast;
  wire        arm_eth1_rx_tready;
  wire [3:0]  arm_eth1_rx_tuser;
  wire [7:0]  arm_eth1_rx_tkeep;

  wire [63:0] arm_eth1_rx_tdata_b;
  wire        arm_eth1_rx_tvalid_b;
  wire        arm_eth1_rx_tlast_b;
  wire        arm_eth1_rx_tready_b;
  wire [3:0]  arm_eth1_rx_tuser_b;
  wire [7:0]  arm_eth1_rx_tkeep_b;

  wire        arm_eth1_tx_irq;
  wire        arm_eth1_rx_irq;

  // Vita to Ethernet
  (* mark_debug ="true" *) wire  [63:0]  v2e0_tdata;
  (* mark_debug ="true" *) wire          v2e0_tlast;
  (* mark_debug ="true" *) wire          v2e0_tvalid;
  (* mark_debug ="true" *) wire          v2e0_tready;

  wire  [63:0]  v2e1_tdata;
  wire          v2e1_tlast;
  wire          v2e1_tvalid;
  wire          v2e1_tready;

  // Ethernet to Vita
  (* mark_debug ="true" *) wire  [63:0]  e2v0_tdata;
  (* mark_debug ="true" *) wire          e2v0_tlast;
  (* mark_debug ="true" *) wire          e2v0_tvalid;
  (* mark_debug ="true" *) wire          e2v0_tready;

  wire  [63:0]  e2v1_tdata;
  wire          e2v1_tlast;
  wire          e2v1_tvalid;
  wire          e2v1_tready;

  /////////////////////////////////////////////////////////////////////
  //
  // Network Interface 0
  //
  //////////////////////////////////////////////////////////////////////

  network_interface #(
`ifdef SFP0_10GBE
      .PROTOCOL("10GbE"),
`elsif SFP0_1GBE
      .PROTOCOL("1GbE"),
`elsif SFP0_AURORA
      .PROTOCOL("Aurora"),
`endif
      .DWIDTH(REG_DWIDTH),     // Width of the AXI4-Lite data bus (must be 32 or 64)
      .AWIDTH(REG_AWIDTH),     // Width of the address bus
      .MDIO_EN(1'b1),
      .PORTNUM(8'd0)
  ) network_interface_0 (
     .areset(global_rst),     // TODO: Add Reset through PS
     .gt_refclk(sfp0_gt_refclk),
     .gb_refclk(sfp0_gb_refclk),
     .misc_clk(sfp0_misc_clk),

     .bus_rst(bus_rst),
     .bus_clk(bus_clk),
   `ifdef SFP0_1GBE
     .gt0_qplloutclk(gt0_qplloutclk),
     .gt0_qplloutrefclk(gt0_qplloutrefclk),
     .pma_reset_out(pma_reset),
   `endif
   `ifdef SFP0_10GBE
     .qplllock(qplllock),
     .qplloutclk(qplloutclk),
     .qplloutrefclk(qplloutrefclk),
   `endif
   `ifdef SFP0_AURORA
     .qplllock(qplllock),
     .qpllreset(qpllreset),
     .qpllrefclklost(qpllrefclklost),
     .qplloutclk(qplloutclk),
     .qplloutrefclk(qplloutrefclk),
   `endif
     .txp(SFP_0_TX_P),
     .txn(SFP_0_TX_N),
     .rxp(SFP_0_RX_P),
     .rxn(SFP_0_RX_N),

     .sfpp_rxlos(SFP_0_LOS),
     .sfpp_tx_fault(SFP_0_TXFAULT),
     .sfpp_tx_disable(SFP_0_TXDISABLE),

     .sfp_phy_status(sfp0_phy_status),

     // Clock and reset
     .s_axi_aclk(clk40),
     .s_axi_aresetn(FCLK_RESET0N),
     // AXI4-Lite: Write address port (domain: s_axi_aclk)
     .s_axi_awaddr(M_AXI_GP0_AWADDR_S1),
     .s_axi_awvalid(M_AXI_GP0_AWVALID_S1),
     .s_axi_awready(M_AXI_GP0_AWREADY_S1),
     // AXI4-Lite: Write data port (domain: s_axi_aclk)
     .s_axi_wdata(M_AXI_GP0_WDATA_S1),
     .s_axi_wstrb(M_AXI_GP0_WSTRB_S1),
     .s_axi_wvalid(M_AXI_GP0_WVALID_S1),
     .s_axi_wready(M_AXI_GP0_WREADY_S1),
     // AXI4-Lite: Write response port (domain: s_axi_aclk)
     .s_axi_bresp(M_AXI_GP0_BRESP_S1),
     .s_axi_bvalid(M_AXI_GP0_BVALID_S1),
     .s_axi_bready(M_AXI_GP0_BREADY_S1),
     // AXI4-Lite: Read address port (domain: s_axi_aclk)
     .s_axi_araddr(M_AXI_GP0_ARADDR_S1),
     .s_axi_arvalid(M_AXI_GP0_ARVALID_S1),
     .s_axi_arready(M_AXI_GP0_ARREADY_S1),
     // AXI4-Lite: Read data port (domain: s_axi_aclk)
     .s_axi_rdata(M_AXI_GP0_RDATA_S1),
     .s_axi_rresp(M_AXI_GP0_RRESP_S1),
     .s_axi_rvalid(M_AXI_GP0_RVALID_S1),
     .s_axi_rready(M_AXI_GP0_RREADY_S1),

     // Ethernet to Vita
     .e2v_tdata(e2v0_tdata),
     .e2v_tlast(e2v0_tlast),
     .e2v_tvalid(e2v0_tvalid),
     .e2v_tready(e2v0_tready),

     // Vita to Ethernet
     .v2e_tdata(v2e0_tdata),
     .v2e_tlast(v2e0_tlast),
     .v2e_tvalid(v2e0_tvalid),
     .v2e_tready(v2e0_tready),

     // Crossover
     .xo_tdata(e01_tdata),
     .xo_tuser(e01_tuser),
     .xo_tlast(e01_tlast),
     .xo_tvalid(e01_tvalid),
     .xo_tready(e01_tready),
     .xi_tdata(e10_tdata),
     .xi_tuser(e10_tuser),
     .xi_tlast(e10_tlast),
     .xi_tvalid(e10_tvalid),
     .xi_tready(e10_tready),

     // Ethernet to CPU
     .e2c_tdata(arm_eth0_rx_tdata_b),
     .e2c_tkeep(arm_eth0_rx_tkeep_b),
     .e2c_tlast(arm_eth0_rx_tlast_b),
     .e2c_tvalid(arm_eth0_rx_tvalid_b),
     .e2c_tready(arm_eth0_rx_tready_b),

     // CPU to Ethernet
     .c2e_tdata(arm_eth0_tx_tdata_b),
     .c2e_tkeep(arm_eth0_tx_tkeep_b),
     .c2e_tlast(arm_eth0_tx_tlast_b),
     .c2e_tvalid(arm_eth0_tx_tvalid_b),
     .c2e_tready(arm_eth0_tx_tready_b),

     // LED
     .activity_led(SFP_0_LED_A)
  );

  /////////////////////////////////////////////////////////////////////
  //
  // Network Interface 1
  //
  //////////////////////////////////////////////////////////////////////

  network_interface #(
`ifdef SFP1_10GBE
      .PROTOCOL("10GbE"),
`elsif SFP1_1GBE
      .PROTOCOL("1GbE"),
`elsif SFP1_AURORA
      .PROTOCOL("Aurora"),
`endif
      .DWIDTH(REG_DWIDTH),     // Width of the AXI4-Lite data bus (must be 32 or 64)
      .AWIDTH(REG_AWIDTH),     // Width of the address bus
      .MDIO_EN(1'b1),
      .PORTNUM(8'd1)
  ) network_interface_1 (
      .areset(global_rst),     // TODO: Add reset through PS
      .gt_refclk(sfp1_gt_refclk),
      .gb_refclk(sfp1_gb_refclk),
      .misc_clk(sfp1_misc_clk),

      .bus_rst(bus_rst),
      .bus_clk(bus_clk),
    `ifdef SFP1_1GBE
      .gt0_qplloutclk(gt0_qplloutclk),
      .gt0_qplloutrefclk(gt0_qplloutrefclk),
      .pma_reset_out(),
    `endif
    `ifdef SFP1_10GBE
      .qpllreset(qpllreset),
      .qplllock(qplllock),
      .qplloutclk(qplloutclk),
      .qplloutrefclk(qplloutrefclk),
    `endif
    `ifdef SFP1_AURORA
      .qplllock(qplllock),
      .qplloutclk(qplloutclk),
      .qplloutrefclk(qplloutrefclk),
     `endif

      .txp(SFP_1_TX_P),
      .txn(SFP_1_TX_N),
      .rxp(SFP_1_RX_P),
      .rxn(SFP_1_RX_N),

      .sfpp_rxlos(SFP_1_LOS),
      .sfpp_tx_fault(SFP_1_TXFAULT),
      .sfpp_tx_disable(SFP_1_TXDISABLE),

      .sfp_phy_status(sfp1_phy_status),

      // Clock and reset
      .s_axi_aclk(clk40),
      .s_axi_aresetn(FCLK_RESET0N),
      // AXI4-Lite: Write address port (domain: s_axi_aclk)
      .s_axi_awaddr(M_AXI_GP0_AWADDR_S3),
      .s_axi_awvalid(M_AXI_GP0_AWVALID_S3),
      .s_axi_awready(M_AXI_GP0_AWREADY_S3),
      // AXI4-Lite: Write data port (domain: s_axi_aclk)
      .s_axi_wdata(M_AXI_GP0_WDATA_S3),
      .s_axi_wstrb(M_AXI_GP0_WSTRB_S3),
      .s_axi_wvalid(M_AXI_GP0_WVALID_S3),
      .s_axi_wready(M_AXI_GP0_WREADY_S3),
      // AXI4-Lite: Write response port (domain: s_axi_aclk)
      .s_axi_bresp(M_AXI_GP0_BRESP_S3),
      .s_axi_bvalid(M_AXI_GP0_BVALID_S3),
      .s_axi_bready(M_AXI_GP0_BREADY_S3),
      // AXI4-Lite: Read address port (domain: s_axi_aclk)
      .s_axi_araddr(M_AXI_GP0_ARADDR_S3),
      .s_axi_arvalid(M_AXI_GP0_ARVALID_S3),
      .s_axi_arready(M_AXI_GP0_ARREADY_S3),
      // AXI4-Lite: Read data port (domain: s_axi_aclk)
      .s_axi_rdata(M_AXI_GP0_RDATA_S3),
      .s_axi_rresp(M_AXI_GP0_RRESP_S3),
      .s_axi_rvalid(M_AXI_GP0_RVALID_S3),
      .s_axi_rready(M_AXI_GP0_RREADY_S3),

      // Ethernet to Vita
      .e2v_tdata(e2v1_tdata),
      .e2v_tlast(e2v1_tlast),
      .e2v_tvalid(e2v1_tvalid),
      .e2v_tready(e2v1_tready),

      // Vita to Ethernet
      .v2e_tdata(v2e1_tdata),
      .v2e_tlast(v2e1_tlast),
      .v2e_tvalid(v2e1_tvalid),
      .v2e_tready(v2e1_tready),

      // Crossover
      .xo_tdata(e10_tdata),
      .xo_tuser(e10_tuser),
      .xo_tlast(e10_tlast),
      .xo_tvalid(e10_tvalid),
      .xo_tready(e10_tready),
      .xi_tdata(e01_tdata),
      .xi_tuser(e01_tuser),
      .xi_tlast(e01_tlast),
      .xi_tvalid(e01_tvalid),
      .xi_tready(e01_tready),

      // Ethernet to CPU
      .e2c_tdata(arm_eth1_rx_tdata_b),
      .e2c_tkeep(arm_eth1_rx_tkeep_b),
      .e2c_tlast(arm_eth1_rx_tlast_b),
      .e2c_tvalid(arm_eth1_rx_tvalid_b),
      .e2c_tready(arm_eth1_rx_tready_b),

      // CPU to Ethernet
      .c2e_tdata(arm_eth1_tx_tdata_b),
      .c2e_tkeep(arm_eth1_tx_tkeep_b),
      .c2e_tlast(arm_eth1_tx_tlast_b),
      .c2e_tvalid(arm_eth1_tx_tvalid_b),
      .c2e_tready(arm_eth1_tx_tready_b),

      // LED
      .activity_led(SFP_1_LED_A)
  );

  /////////////////////////////////////////////////////////////////////
  //
  // Ethernet DMA 0
  //
  //////////////////////////////////////////////////////////////////////

  assign  IRQ_F2P[0] = arm_eth0_rx_irq;
  assign  IRQ_F2P[1] = arm_eth0_tx_irq;

  assign {S_AXI_HP0_AWID, S_AXI_HP0_ARID} = 12'd0;
  assign {S_AXI_GP0_AWID, S_AXI_GP0_ARID} = 12'd0;

  axi_eth_dma inst_axi_eth_dma0
  (
    .s_axi_lite_aclk(clk40),
    .m_axi_sg_aclk(clk40),
    .m_axi_mm2s_aclk(clk40),
    .m_axi_s2mm_aclk(clk40),
    .axi_resetn(FCLK_RESET0N),

    .s_axi_lite_awaddr(M_AXI_GP0_AWADDR_S0),
    .s_axi_lite_awvalid(M_AXI_GP0_AWVALID_S0),
    .s_axi_lite_awready(M_AXI_GP0_AWREADY_S0),

    .s_axi_lite_wdata(M_AXI_GP0_WDATA_S0),
    .s_axi_lite_wvalid(M_AXI_GP0_WVALID_S0),
    .s_axi_lite_wready(M_AXI_GP0_WREADY_S0),

    .s_axi_lite_bresp(M_AXI_GP0_BRESP_S0),
    .s_axi_lite_bvalid(M_AXI_GP0_BVALID_S0),
    .s_axi_lite_bready(M_AXI_GP0_BREADY_S0),

    .s_axi_lite_araddr(M_AXI_GP0_ARADDR_S0),
    .s_axi_lite_arvalid(M_AXI_GP0_ARVALID_S0),
    .s_axi_lite_arready(M_AXI_GP0_ARREADY_S0),

    .s_axi_lite_rdata(M_AXI_GP0_RDATA_S0),
    .s_axi_lite_rresp(M_AXI_GP0_RRESP_S0),
    .s_axi_lite_rvalid(M_AXI_GP0_RVALID_S0),
    .s_axi_lite_rready(M_AXI_GP0_RREADY_S0),

    .m_axi_sg_awaddr(S_AXI_GP0_AWADDR),
    .m_axi_sg_awlen(S_AXI_GP0_AWLEN),
    .m_axi_sg_awsize(S_AXI_GP0_AWSIZE),
    .m_axi_sg_awburst(S_AXI_GP0_AWBURST),
    .m_axi_sg_awprot(S_AXI_GP0_AWPROT),
    .m_axi_sg_awcache(S_AXI_GP0_AWCACHE),
    .m_axi_sg_awvalid(S_AXI_GP0_AWVALID),
    .m_axi_sg_awready(S_AXI_GP0_AWREADY),
    .m_axi_sg_wdata(S_AXI_GP0_WDATA),
    .m_axi_sg_wstrb(S_AXI_GP0_WSTRB),
    .m_axi_sg_wlast(S_AXI_GP0_WLAST),
    .m_axi_sg_wvalid(S_AXI_GP0_WVALID),
    .m_axi_sg_wready(S_AXI_GP0_WREADY),
    .m_axi_sg_bresp(S_AXI_GP0_BRESP),
    .m_axi_sg_bvalid(S_AXI_GP0_BVALID),
    .m_axi_sg_bready(S_AXI_GP0_BREADY),
    .m_axi_sg_araddr(S_AXI_GP0_ARADDR),
    .m_axi_sg_arlen(S_AXI_GP0_ARLEN),
    .m_axi_sg_arsize(S_AXI_GP0_ARSIZE),
    .m_axi_sg_arburst(S_AXI_GP0_ARBURST),
    .m_axi_sg_arprot(S_AXI_GP0_ARPROT),
    .m_axi_sg_arcache(S_AXI_GP0_ARCACHE),
    .m_axi_sg_arvalid(S_AXI_GP0_ARVALID),
    .m_axi_sg_arready(S_AXI_GP0_ARREADY),
    .m_axi_sg_rdata(S_AXI_GP0_RDATA),
    .m_axi_sg_rresp(S_AXI_GP0_RRESP),
    .m_axi_sg_rlast(S_AXI_GP0_RLAST),
    .m_axi_sg_rvalid(S_AXI_GP0_RVALID),
    .m_axi_sg_rready(S_AXI_GP0_RREADY),

    .m_axi_mm2s_araddr(S_AXI_HP0_ARADDR),
    .m_axi_mm2s_arlen(S_AXI_HP0_ARLEN),
    .m_axi_mm2s_arsize(S_AXI_HP0_ARSIZE),
    .m_axi_mm2s_arburst(S_AXI_HP0_ARBURST),
    .m_axi_mm2s_arprot(S_AXI_HP0_ARPROT),
    .m_axi_mm2s_arcache(S_AXI_HP0_ARCACHE),
    .m_axi_mm2s_arvalid(S_AXI_HP0_ARVALID),
    .m_axi_mm2s_arready(S_AXI_HP0_ARREADY),
    .m_axi_mm2s_rdata(S_AXI_HP0_RDATA),
    .m_axi_mm2s_rresp(S_AXI_HP0_RRESP),
    .m_axi_mm2s_rlast(S_AXI_HP0_RLAST),
    .m_axi_mm2s_rvalid(S_AXI_HP0_RVALID),
    .m_axi_mm2s_rready(S_AXI_HP0_RREADY),

    .mm2s_prmry_reset_out_n(),
    .m_axis_mm2s_tdata(arm_eth0_tx_tdata),
    .m_axis_mm2s_tkeep(arm_eth0_tx_tkeep),
    .m_axis_mm2s_tvalid(arm_eth0_tx_tvalid),
    .m_axis_mm2s_tready(arm_eth0_tx_tready),
    .m_axis_mm2s_tlast(arm_eth0_tx_tlast),

    .m_axi_s2mm_awaddr(S_AXI_HP0_AWADDR),
    .m_axi_s2mm_awlen(S_AXI_HP0_AWLEN),
    .m_axi_s2mm_awsize(S_AXI_HP0_AWSIZE),
    .m_axi_s2mm_awburst(S_AXI_HP0_AWBURST),
    .m_axi_s2mm_awprot(S_AXI_HP0_AWPROT),
    .m_axi_s2mm_awcache(S_AXI_HP0_AWCACHE),
    .m_axi_s2mm_awvalid(S_AXI_HP0_AWVALID),
    .m_axi_s2mm_awready(S_AXI_HP0_AWREADY),
    .m_axi_s2mm_wdata(S_AXI_HP0_WDATA),
    .m_axi_s2mm_wstrb(S_AXI_HP0_WSTRB),
    .m_axi_s2mm_wlast(S_AXI_HP0_WLAST),
    .m_axi_s2mm_wvalid(S_AXI_HP0_WVALID),
    .m_axi_s2mm_wready(S_AXI_HP0_WREADY),
    .m_axi_s2mm_bresp(S_AXI_HP0_BRESP),
    .m_axi_s2mm_bvalid(S_AXI_HP0_BVALID),
    .m_axi_s2mm_bready(S_AXI_HP0_BREADY),

    .s2mm_prmry_reset_out_n(),
    .s_axis_s2mm_tdata(arm_eth0_rx_tdata),
    .s_axis_s2mm_tkeep(arm_eth0_rx_tkeep),
    .s_axis_s2mm_tvalid(arm_eth0_rx_tvalid),
    .s_axis_s2mm_tready(arm_eth0_rx_tready),
    .s_axis_s2mm_tlast(arm_eth0_rx_tlast),

    .mm2s_introut(arm_eth0_tx_irq),
    .s2mm_introut(arm_eth0_rx_irq),
    .axi_dma_tstvec()
  );

  axis_fifo_2clk #( .WIDTH(1+8+64)) eth_tx_0_fifo_2clk_i (
    .s_axis_areset(FCLK_RESET0), .s_axis_aclk(clk40),
    .s_axis_tdata({arm_eth0_tx_tlast, arm_eth0_tx_tkeep, arm_eth0_tx_tdata}),
    .s_axis_tvalid(arm_eth0_tx_tvalid),
    .s_axis_tready(arm_eth0_tx_tready),
    .m_axis_aclk(bus_clk),
    .m_axis_tdata({arm_eth0_tx_tlast_b, arm_eth0_tx_tkeep_b, arm_eth0_tx_tdata_b}),
    .m_axis_tvalid(arm_eth0_tx_tvalid_b),
    .m_axis_tready(arm_eth0_tx_tready_b)
  );

  axis_fifo_2clk #( .WIDTH(1+8+64)) eth_rx_0_fifo_2clk_i (
    .s_axis_areset(bus_rst), .s_axis_aclk(bus_clk),
    .s_axis_tdata({arm_eth0_rx_tlast_b, arm_eth0_rx_tkeep_b, arm_eth0_rx_tdata_b}),
    .s_axis_tvalid(arm_eth0_rx_tvalid_b),
    .s_axis_tready(arm_eth0_rx_tready_b),
    .m_axis_aclk(clk40),
    .m_axis_tdata({arm_eth0_rx_tlast, arm_eth0_rx_tkeep, arm_eth0_rx_tdata}),
    .m_axis_tvalid(arm_eth0_rx_tvalid),
    .m_axis_tready(arm_eth0_rx_tready)
  );

  /////////////////////////////////////////////////////////////////////
  //
  // Ethernet DMA 1
  //
  //////////////////////////////////////////////////////////////////////

  assign  IRQ_F2P[2] = arm_eth1_rx_irq;
  assign  IRQ_F2P[3] = arm_eth1_tx_irq;

  assign {S_AXI_HP1_AWID, S_AXI_HP1_ARID} = 12'd0;
  assign {S_AXI_GP1_AWID, S_AXI_GP1_ARID} = 12'd0;

  axi_eth_dma inst_axi_eth_dma1
  (
    .s_axi_lite_aclk(clk40),
    .m_axi_sg_aclk(clk40),
    .m_axi_mm2s_aclk(clk40),
    .m_axi_s2mm_aclk(clk40),
    .axi_resetn(FCLK_RESET0N),

    .s_axi_lite_awaddr(M_AXI_GP0_AWADDR_S2),
    .s_axi_lite_awvalid(M_AXI_GP0_AWVALID_S2),
    .s_axi_lite_awready(M_AXI_GP0_AWREADY_S2),

    .s_axi_lite_wdata(M_AXI_GP0_WDATA_S2),
    .s_axi_lite_wvalid(M_AXI_GP0_WVALID_S2),
    .s_axi_lite_wready(M_AXI_GP0_WREADY_S2),

    .s_axi_lite_bresp(M_AXI_GP0_BRESP_S2),
    .s_axi_lite_bvalid(M_AXI_GP0_BVALID_S2),
    .s_axi_lite_bready(M_AXI_GP0_BREADY_S2),

    .s_axi_lite_araddr(M_AXI_GP0_ARADDR_S2),
    .s_axi_lite_arvalid(M_AXI_GP0_ARVALID_S2),
    .s_axi_lite_arready(M_AXI_GP0_ARREADY_S2),

    .s_axi_lite_rdata(M_AXI_GP0_RDATA_S2),
    .s_axi_lite_rresp(M_AXI_GP0_RRESP_S2),
    .s_axi_lite_rvalid(M_AXI_GP0_RVALID_S2),
    .s_axi_lite_rready(M_AXI_GP0_RREADY_S2),

    .m_axi_sg_awaddr(S_AXI_GP1_AWADDR),
    .m_axi_sg_awlen(S_AXI_GP1_AWLEN),
    .m_axi_sg_awsize(S_AXI_GP1_AWSIZE),
    .m_axi_sg_awburst(S_AXI_GP1_AWBURST),
    .m_axi_sg_awprot(S_AXI_GP1_AWPROT),
    .m_axi_sg_awcache(S_AXI_GP1_AWCACHE),
    .m_axi_sg_awvalid(S_AXI_GP1_AWVALID),
    .m_axi_sg_awready(S_AXI_GP1_AWREADY),
    .m_axi_sg_wdata(S_AXI_GP1_WDATA),
    .m_axi_sg_wstrb(S_AXI_GP1_WSTRB),
    .m_axi_sg_wlast(S_AXI_GP1_WLAST),
    .m_axi_sg_wvalid(S_AXI_GP1_WVALID),
    .m_axi_sg_wready(S_AXI_GP1_WREADY),
    .m_axi_sg_bresp(S_AXI_GP1_BRESP),
    .m_axi_sg_bvalid(S_AXI_GP1_BVALID),
    .m_axi_sg_bready(S_AXI_GP1_BREADY),
    .m_axi_sg_araddr(S_AXI_GP1_ARADDR),
    .m_axi_sg_arlen(S_AXI_GP1_ARLEN),
    .m_axi_sg_arsize(S_AXI_GP1_ARSIZE),
    .m_axi_sg_arburst(S_AXI_GP1_ARBURST),
    .m_axi_sg_arprot(S_AXI_GP1_ARPROT),
    .m_axi_sg_arcache(S_AXI_GP1_ARCACHE),
    .m_axi_sg_arvalid(S_AXI_GP1_ARVALID),
    .m_axi_sg_arready(S_AXI_GP1_ARREADY),
    .m_axi_sg_rdata(S_AXI_GP1_RDATA),
    .m_axi_sg_rresp(S_AXI_GP1_RRESP),
    .m_axi_sg_rlast(S_AXI_GP1_RLAST),
    .m_axi_sg_rvalid(S_AXI_GP1_RVALID),
    .m_axi_sg_rready(S_AXI_GP1_RREADY),

    .m_axi_mm2s_araddr(S_AXI_HP1_ARADDR),
    .m_axi_mm2s_arlen(S_AXI_HP1_ARLEN),
    .m_axi_mm2s_arsize(S_AXI_HP1_ARSIZE),
    .m_axi_mm2s_arburst(S_AXI_HP1_ARBURST),
    .m_axi_mm2s_arprot(S_AXI_HP1_ARPROT),
    .m_axi_mm2s_arcache(S_AXI_HP1_ARCACHE),
    .m_axi_mm2s_arvalid(S_AXI_HP1_ARVALID),
    .m_axi_mm2s_arready(S_AXI_HP1_ARREADY),
    .m_axi_mm2s_rdata(S_AXI_HP1_RDATA),
    .m_axi_mm2s_rresp(S_AXI_HP1_RRESP),
    .m_axi_mm2s_rlast(S_AXI_HP1_RLAST),
    .m_axi_mm2s_rvalid(S_AXI_HP1_RVALID),
    .m_axi_mm2s_rready(S_AXI_HP1_RREADY),

    .mm2s_prmry_reset_out_n(),
    .m_axis_mm2s_tdata(arm_eth1_tx_tdata),
    .m_axis_mm2s_tkeep(arm_eth1_tx_tkeep),
    .m_axis_mm2s_tvalid(arm_eth1_tx_tvalid),
    .m_axis_mm2s_tready(arm_eth1_tx_tready),
    .m_axis_mm2s_tlast(arm_eth1_tx_tlast),

    .m_axi_s2mm_awaddr(S_AXI_HP1_AWADDR),
    .m_axi_s2mm_awlen(S_AXI_HP1_AWLEN),
    .m_axi_s2mm_awsize(S_AXI_HP1_AWSIZE),
    .m_axi_s2mm_awburst(S_AXI_HP1_AWBURST),
    .m_axi_s2mm_awprot(S_AXI_HP1_AWPROT),
    .m_axi_s2mm_awcache(S_AXI_HP1_AWCACHE),
    .m_axi_s2mm_awvalid(S_AXI_HP1_AWVALID),
    .m_axi_s2mm_awready(S_AXI_HP1_AWREADY),
    .m_axi_s2mm_wdata(S_AXI_HP1_WDATA),
    .m_axi_s2mm_wstrb(S_AXI_HP1_WSTRB),
    .m_axi_s2mm_wlast(S_AXI_HP1_WLAST),
    .m_axi_s2mm_wvalid(S_AXI_HP1_WVALID),
    .m_axi_s2mm_wready(S_AXI_HP1_WREADY),
    .m_axi_s2mm_bresp(S_AXI_HP1_BRESP),
    .m_axi_s2mm_bvalid(S_AXI_HP1_BVALID),
    .m_axi_s2mm_bready(S_AXI_HP1_BREADY),

    .s2mm_prmry_reset_out_n(),
    .s_axis_s2mm_tdata(arm_eth1_rx_tdata),
    .s_axis_s2mm_tkeep(arm_eth1_rx_tkeep),
    .s_axis_s2mm_tvalid(arm_eth1_rx_tvalid),
    .s_axis_s2mm_tready(arm_eth1_rx_tready),
    .s_axis_s2mm_tlast(arm_eth1_rx_tlast),

    .mm2s_introut(arm_eth1_tx_irq),
    .s2mm_introut(arm_eth1_rx_irq),
    .axi_dma_tstvec()
  );

  axis_fifo_2clk #( .WIDTH(1+8+64)) eth_tx_1_fifo_2clk_i (
    .s_axis_areset(FCLK_RESET0), .s_axis_aclk(clk40),
    .s_axis_tdata({arm_eth1_tx_tlast, arm_eth1_tx_tkeep, arm_eth1_tx_tdata}),
    .s_axis_tvalid(arm_eth1_tx_tvalid),
    .s_axis_tready(arm_eth1_tx_tready),
    .m_axis_aclk(bus_clk),
    .m_axis_tdata({arm_eth1_tx_tlast_b, arm_eth1_tx_tkeep_b, arm_eth1_tx_tdata_b}),
    .m_axis_tvalid(arm_eth1_tx_tvalid_b),
    .m_axis_tready(arm_eth1_tx_tready_b)
  );

  axis_fifo_2clk #( .WIDTH(1+8+64)) eth_rx_1_fifo_2clk_i (
    .s_axis_areset(bus_rst), .s_axis_aclk(bus_clk),
    .s_axis_tdata({arm_eth1_rx_tlast_b, arm_eth1_rx_tkeep_b, arm_eth1_rx_tdata_b}),
    .s_axis_tvalid(arm_eth1_rx_tvalid_b),
    .s_axis_tready(arm_eth1_rx_tready_b),
    .m_axis_aclk(clk40),
    .m_axis_tdata({arm_eth1_rx_tlast, arm_eth1_rx_tkeep, arm_eth1_rx_tdata}),
    .m_axis_tvalid(arm_eth1_rx_tvalid),
    .m_axis_tready(arm_eth1_rx_tready)
  );

  /////////////////////////////////////////////////////////////////////
  //
  // AXI Interconnect
  //
  // Slave 0: Ethernet DMA 0
  // Slave 1: Network Interface 0
  // Slave 2: Ethernet DMA 1
  // Slave 3: Network Interface 1
  // Slave 4: XBAR
  // Slave 5: Clocking and Jesd Core
  // Slave 6: XBAR DMA
  //
  //////////////////////////////////////////////////////////////////////

  axi_interconnect inst_axi_interconnect
  (
    .aclk(clk40),
    .aresetn(FCLK_RESET0N),
    .s_axi_awaddr(M_AXI_GP0_AWADDR),
    .s_axi_awprot(3'b0),               //Recommended default value
    .s_axi_awready(M_AXI_GP0_AWREADY),
    .s_axi_awvalid(M_AXI_GP0_AWVALID),
    .s_axi_wdata(M_AXI_GP0_WDATA),
    .s_axi_wstrb(M_AXI_GP0_WSTRB),
    .s_axi_wvalid(M_AXI_GP0_WVALID),
    .s_axi_wready(M_AXI_GP0_WREADY),
    .s_axi_bresp(M_AXI_GP0_BRESP),
    .s_axi_bvalid(M_AXI_GP0_BVALID),
    .s_axi_bready(M_AXI_GP0_BREADY),
    .s_axi_araddr(M_AXI_GP0_ARADDR),
    .s_axi_arprot(3'b0),               //Recommended default value
    .s_axi_arvalid(M_AXI_GP0_ARVALID),
    .s_axi_arready(M_AXI_GP0_ARREADY),
    .s_axi_rdata(M_AXI_GP0_RDATA),
    .s_axi_rresp(M_AXI_GP0_RRESP),
    .s_axi_rvalid(M_AXI_GP0_RVALID),
    .s_axi_rready(M_AXI_GP0_RREADY),
    .m_axi_awaddr({M_AXI_GP0_AWADDR_S6, M_AXI_GP0_AWADDR_S5, M_AXI_GP0_AWADDR_S4, M_AXI_GP0_AWADDR_S3, M_AXI_GP0_AWADDR_S2, M_AXI_GP0_AWADDR_S1, M_AXI_GP0_AWADDR_S0}),
    .m_axi_awvalid({M_AXI_GP0_AWVALID_S6, M_AXI_GP0_AWVALID_S5, M_AXI_GP0_AWVALID_S4, M_AXI_GP0_AWVALID_S3, M_AXI_GP0_AWVALID_S2, M_AXI_GP0_AWVALID_S1, M_AXI_GP0_AWVALID_S0}),
    .m_axi_awready({M_AXI_GP0_AWREADY_S6, M_AXI_GP0_AWREADY_S5, M_AXI_GP0_AWREADY_S4, M_AXI_GP0_AWREADY_S3, M_AXI_GP0_AWREADY_S2, M_AXI_GP0_AWREADY_S1, M_AXI_GP0_AWREADY_S0}),
    .m_axi_wdata({M_AXI_GP0_WDATA_S6, M_AXI_GP0_WDATA_S5, M_AXI_GP0_WDATA_S4, M_AXI_GP0_WDATA_S3, M_AXI_GP0_WDATA_S2, M_AXI_GP0_WDATA_S1, M_AXI_GP0_WDATA_S0}),
    .m_axi_wstrb({M_AXI_GP0_WSTRB_S6, M_AXI_GP0_WSTRB_S5, M_AXI_GP0_WSTRB_S4, M_AXI_GP0_WSTRB_S3, M_AXI_GP0_WSTRB_S2, M_AXI_GP0_WSTRB_S1, M_AXI_GP0_WSTRB_S0}),
    .m_axi_wvalid({M_AXI_GP0_WVALID_S6, M_AXI_GP0_WVALID_S5, M_AXI_GP0_WVALID_S4, M_AXI_GP0_WVALID_S3, M_AXI_GP0_WVALID_S2, M_AXI_GP0_WVALID_S1, M_AXI_GP0_WVALID_S0}),
    .m_axi_wready({M_AXI_GP0_WREADY_S6, M_AXI_GP0_WREADY_S5, M_AXI_GP0_WREADY_S4, M_AXI_GP0_WREADY_S3, M_AXI_GP0_WREADY_S2, M_AXI_GP0_WREADY_S1, M_AXI_GP0_WREADY_S0}),
    .m_axi_bresp({M_AXI_GP0_BRESP_S6, M_AXI_GP0_BRESP_S5, M_AXI_GP0_BRESP_S4, M_AXI_GP0_BRESP_S3, M_AXI_GP0_BRESP_S2, M_AXI_GP0_BRESP_S1, M_AXI_GP0_BRESP_S0}),
    .m_axi_bvalid({M_AXI_GP0_BVALID_S6, M_AXI_GP0_BVALID_S5, M_AXI_GP0_BVALID_S4, M_AXI_GP0_BVALID_S3, M_AXI_GP0_BVALID_S2, M_AXI_GP0_BVALID_S1, M_AXI_GP0_BVALID_S0}),
    .m_axi_bready({M_AXI_GP0_BREADY_S6, M_AXI_GP0_BREADY_S5, M_AXI_GP0_BREADY_S4, M_AXI_GP0_BREADY_S3, M_AXI_GP0_BREADY_S2, M_AXI_GP0_BREADY_S1, M_AXI_GP0_BREADY_S0}),
    .m_axi_araddr({M_AXI_GP0_ARADDR_S6, M_AXI_GP0_ARADDR_S5, M_AXI_GP0_ARADDR_S4, M_AXI_GP0_ARADDR_S3, M_AXI_GP0_ARADDR_S2, M_AXI_GP0_ARADDR_S1, M_AXI_GP0_ARADDR_S0}),
    .m_axi_arvalid({M_AXI_GP0_ARVALID_S6, M_AXI_GP0_ARVALID_S5, M_AXI_GP0_ARVALID_S4, M_AXI_GP0_ARVALID_S3, M_AXI_GP0_ARVALID_S2, M_AXI_GP0_ARVALID_S1, M_AXI_GP0_ARVALID_S0}),
    .m_axi_arready({M_AXI_GP0_ARREADY_S6, M_AXI_GP0_ARREADY_S5, M_AXI_GP0_ARREADY_S4, M_AXI_GP0_ARREADY_S3, M_AXI_GP0_ARREADY_S2, M_AXI_GP0_ARREADY_S1, M_AXI_GP0_ARREADY_S0}),
    .m_axi_rdata({M_AXI_GP0_RDATA_S6, M_AXI_GP0_RDATA_S5, M_AXI_GP0_RDATA_S4, M_AXI_GP0_RDATA_S3, M_AXI_GP0_RDATA_S2, M_AXI_GP0_RDATA_S1, M_AXI_GP0_RDATA_S0}),
    .m_axi_rresp({M_AXI_GP0_RRESP_S6, M_AXI_GP0_RRESP_S5, M_AXI_GP0_RRESP_S4, M_AXI_GP0_RRESP_S3, M_AXI_GP0_RRESP_S2, M_AXI_GP0_RRESP_S1, M_AXI_GP0_RRESP_S0}),
    .m_axi_rvalid({M_AXI_GP0_RVALID_S6, M_AXI_GP0_RVALID_S5, M_AXI_GP0_RVALID_S4, M_AXI_GP0_RVALID_S3, M_AXI_GP0_RVALID_S2, M_AXI_GP0_RVALID_S1, M_AXI_GP0_RVALID_S0}),
    .m_axi_rready({M_AXI_GP0_RREADY_S6, M_AXI_GP0_RREADY_S5, M_AXI_GP0_RREADY_S4, M_AXI_GP0_RREADY_S3, M_AXI_GP0_RREADY_S2, M_AXI_GP0_RREADY_S1, M_AXI_GP0_RREADY_S0})
  );

  /////////////////////////////////////////////////////////////////////
  //
  // Processing System
  //
  //////////////////////////////////////////////////////////////////////

  wire spi0_sclk;
  wire spi0_mosi;
  wire spi0_miso;
  wire spi0_ss0;
  wire spi0_ss1;
  wire spi0_ss2;
  wire spi1_sclk;
  wire spi1_mosi;
  wire spi1_miso;
  wire spi1_ss0;
  wire spi1_ss1;
  wire spi1_ss2;

  wire [63:0] ps_gpio_out;
  wire [63:0] ps_gpio_in;
  wire [63:0] ps_gpio_tri;

  assign DBA_CPLD_JTAG_TCK = ps_gpio_out[0];
  assign DBA_CPLD_JTAG_TDI = ps_gpio_out[1];
  assign DBA_CPLD_JTAG_TMS = ps_gpio_out[2];
  assign ps_gpio_in[3]     = DBA_CPLD_JTAG_TDO;

  assign DBB_CPLD_JTAG_TCK = ps_gpio_out[4];
  assign DBB_CPLD_JTAG_TDI = ps_gpio_out[5];
  assign DBB_CPLD_JTAG_TMS = ps_gpio_out[6];
  assign ps_gpio_in[7]     = DBB_CPLD_JTAG_TDO;

  genvar i;
  generate for (i=0; i<12; i=i+1) begin: io_tristate_gen
    assign FPGA_GPIO[i] = ps_gpio_tri[32+i] ? 1'bz : ps_gpio_out[32+i];
    assign ps_gpio_in[32+i] = FPGA_GPIO[i];
  end endgenerate

  n310_ps inst_n310_ps
  (
    .SPI0_SCLK(spi0_sclk),
    .SPI0_MOSI(spi0_mosi),
    .SPI0_MISO(spi0_miso),
    .SPI0_SS0(spi0_ss0),
    .SPI0_SS1(spi0_ss1),
    .SPI0_SS2(spi0_ss2),

    .SPI1_SCLK(spi1_sclk),
    .SPI1_MOSI(spi1_mosi),
    .SPI1_MISO(spi1_miso),
    .SPI1_SS0(spi1_ss0),
    .SPI1_SS1(spi1_ss1),
    .SPI1_SS2(spi1_ss2),

    .M_AXI_GP0_ARVALID(M_AXI_GP0_ARVALID),
    .M_AXI_GP0_ARREADY(M_AXI_GP0_ARREADY),
    .M_AXI_GP0_ARADDR(M_AXI_GP0_ARADDR),
     // Write Address Channel
    .M_AXI_GP0_AWVALID(M_AXI_GP0_AWVALID),
    .M_AXI_GP0_AWREADY(M_AXI_GP0_AWREADY),
    .M_AXI_GP0_AWADDR(M_AXI_GP0_AWADDR),
    // Write Data Channel
    .M_AXI_GP0_WVALID(M_AXI_GP0_WVALID),
    .M_AXI_GP0_WDATA(M_AXI_GP0_WDATA),
    .M_AXI_GP0_WSTRB(M_AXI_GP0_WSTRB),
    .M_AXI_GP0_WREADY(M_AXI_GP0_WREADY),
    // Read Data Channel
    .M_AXI_GP0_RVALID(M_AXI_GP0_RVALID),
    .M_AXI_GP0_RDATA(M_AXI_GP0_RDATA),
    .M_AXI_GP0_RRESP(M_AXI_GP0_RRESP),
    .M_AXI_GP0_RREADY(M_AXI_GP0_RREADY),
    // Write Response Channel
    .M_AXI_GP0_BREADY(M_AXI_GP0_BREADY),
    .M_AXI_GP0_BRESP(M_AXI_GP0_BRESP),
    .M_AXI_GP0_BVALID(M_AXI_GP0_BVALID),

    .S_AXI_HP0_AWID(S_AXI_HP0_AWID),
    .S_AXI_HP0_AWADDR(S_AXI_HP0_AWADDR),
    .S_AXI_HP0_AWPROT(S_AXI_HP0_AWPROT),
    .S_AXI_HP0_AWVALID(S_AXI_HP0_AWVALID),
    .S_AXI_HP0_AWREADY(S_AXI_HP0_AWREADY),
    .S_AXI_HP0_WDATA(S_AXI_HP0_WDATA),
    .S_AXI_HP0_WSTRB(S_AXI_HP0_WSTRB),
    .S_AXI_HP0_WVALID(S_AXI_HP0_WVALID),
    .S_AXI_HP0_WREADY(S_AXI_HP0_WREADY),
    .S_AXI_HP0_BRESP(S_AXI_HP0_BRESP),
    .S_AXI_HP0_BVALID(S_AXI_HP0_BVALID),
    .S_AXI_HP0_BREADY(S_AXI_HP0_BREADY),
    .S_AXI_HP0_ARID(S_AXI_HP0_ARID),
    .S_AXI_HP0_ARADDR(S_AXI_HP0_ARADDR),
    .S_AXI_HP0_ARPROT(S_AXI_HP0_ARPROT),
    .S_AXI_HP0_ARVALID(S_AXI_HP0_ARVALID),
    .S_AXI_HP0_ARREADY(S_AXI_HP0_ARREADY),
    .S_AXI_HP0_RDATA(S_AXI_HP0_RDATA),
    .S_AXI_HP0_RRESP(S_AXI_HP0_RRESP),
    .S_AXI_HP0_RVALID(S_AXI_HP0_RVALID),
    .S_AXI_HP0_RREADY(S_AXI_HP0_RREADY),
    .S_AXI_HP0_AWLEN(S_AXI_HP0_AWLEN),
    .S_AXI_HP0_RLAST(S_AXI_HP0_RLAST),
    .S_AXI_HP0_ARCACHE(S_AXI_HP0_ARCACHE),
    .S_AXI_HP0_AWSIZE(S_AXI_HP0_AWSIZE),
    .S_AXI_HP0_AWBURST(S_AXI_HP0_AWBURST),
    .S_AXI_HP0_AWCACHE(S_AXI_HP0_AWCACHE),
    .S_AXI_HP0_WLAST(S_AXI_HP0_WLAST),
    .S_AXI_HP0_ARLEN(S_AXI_HP0_ARLEN),
    .S_AXI_HP0_ARBURST(S_AXI_HP0_ARBURST),
    .S_AXI_HP0_ARSIZE(S_AXI_HP0_ARSIZE),

    .S_AXI_GP0_AWID(S_AXI_GP0_AWID),
    .S_AXI_GP0_AWADDR(S_AXI_GP0_AWADDR),
    .S_AXI_GP0_AWPROT(S_AXI_GP0_AWPROT),
    .S_AXI_GP0_AWVALID(S_AXI_GP0_AWVALID),
    .S_AXI_GP0_AWREADY(S_AXI_GP0_AWREADY),
    .S_AXI_GP0_WDATA(S_AXI_GP0_WDATA),
    .S_AXI_GP0_WSTRB(S_AXI_GP0_WSTRB),
    .S_AXI_GP0_WVALID(S_AXI_GP0_WVALID),
    .S_AXI_GP0_WREADY(S_AXI_GP0_WREADY),
    .S_AXI_GP0_BRESP(S_AXI_GP0_BRESP),
    .S_AXI_GP0_BVALID(S_AXI_GP0_BVALID),
    .S_AXI_GP0_BREADY(S_AXI_GP0_BREADY),
    .S_AXI_GP0_ARID(S_AXI_GP0_ARID),
    .S_AXI_GP0_ARADDR(S_AXI_GP0_ARADDR),
    .S_AXI_GP0_ARPROT(S_AXI_GP0_ARPROT),
    .S_AXI_GP0_ARVALID(S_AXI_GP0_ARVALID),
    .S_AXI_GP0_ARREADY(S_AXI_GP0_ARREADY),
    .S_AXI_GP0_RDATA(S_AXI_GP0_RDATA),
    .S_AXI_GP0_RRESP(S_AXI_GP0_RRESP),
    .S_AXI_GP0_RVALID(S_AXI_GP0_RVALID),
    .S_AXI_GP0_RREADY(S_AXI_GP0_RREADY),
    .S_AXI_GP0_AWLEN(S_AXI_GP0_AWLEN),
    .S_AXI_GP0_RLAST(S_AXI_GP0_RLAST),
    .S_AXI_GP0_ARCACHE(S_AXI_GP0_ARCACHE),
    .S_AXI_GP0_AWSIZE(S_AXI_GP0_AWSIZE),
    .S_AXI_GP0_AWBURST(S_AXI_GP0_AWBURST),
    .S_AXI_GP0_AWCACHE(S_AXI_GP0_AWCACHE),
    .S_AXI_GP0_WLAST(S_AXI_GP0_WLAST),
    .S_AXI_GP0_ARLEN(S_AXI_GP0_ARLEN),
    .S_AXI_GP0_ARBURST(S_AXI_GP0_ARBURST),
    .S_AXI_GP0_ARSIZE(S_AXI_GP0_ARSIZE),

    .S_AXI_HP1_AWID(S_AXI_HP1_AWID),
    .S_AXI_HP1_AWADDR(S_AXI_HP1_AWADDR),
    .S_AXI_HP1_AWPROT(S_AXI_HP1_AWPROT),
    .S_AXI_HP1_AWVALID(S_AXI_HP1_AWVALID),
    .S_AXI_HP1_AWREADY(S_AXI_HP1_AWREADY),
    .S_AXI_HP1_WDATA(S_AXI_HP1_WDATA),
    .S_AXI_HP1_WSTRB(S_AXI_HP1_WSTRB),
    .S_AXI_HP1_WVALID(S_AXI_HP1_WVALID),
    .S_AXI_HP1_WREADY(S_AXI_HP1_WREADY),
    .S_AXI_HP1_BRESP(S_AXI_HP1_BRESP),
    .S_AXI_HP1_BVALID(S_AXI_HP1_BVALID),
    .S_AXI_HP1_BREADY(S_AXI_HP1_BREADY),
    .S_AXI_HP1_ARID(S_AXI_HP1_ARID),
    .S_AXI_HP1_ARADDR(S_AXI_HP1_ARADDR),
    .S_AXI_HP1_ARPROT(S_AXI_HP1_ARPROT),
    .S_AXI_HP1_ARVALID(S_AXI_HP1_ARVALID),
    .S_AXI_HP1_ARREADY(S_AXI_HP1_ARREADY),
    .S_AXI_HP1_RDATA(S_AXI_HP1_RDATA),
    .S_AXI_HP1_RRESP(S_AXI_HP1_RRESP),
    .S_AXI_HP1_RVALID(S_AXI_HP1_RVALID),
    .S_AXI_HP1_RREADY(S_AXI_HP1_RREADY),
    .S_AXI_HP1_AWLEN(S_AXI_HP1_AWLEN),
    .S_AXI_HP1_RLAST(S_AXI_HP1_RLAST),
    .S_AXI_HP1_ARCACHE(S_AXI_HP1_ARCACHE),
    .S_AXI_HP1_AWSIZE(S_AXI_HP1_AWSIZE),
    .S_AXI_HP1_AWBURST(S_AXI_HP1_AWBURST),
    .S_AXI_HP1_AWCACHE(S_AXI_HP1_AWCACHE),
    .S_AXI_HP1_WLAST(S_AXI_HP1_WLAST),
    .S_AXI_HP1_ARLEN(S_AXI_HP1_ARLEN),
    .S_AXI_HP1_ARBURST(S_AXI_HP1_ARBURST),
    .S_AXI_HP1_ARSIZE(S_AXI_HP1_ARSIZE),

    .S_AXI_GP1_AWID(S_AXI_GP1_AWID),
    .S_AXI_GP1_AWADDR(S_AXI_GP1_AWADDR),
    .S_AXI_GP1_AWPROT(S_AXI_GP1_AWPROT),
    .S_AXI_GP1_AWVALID(S_AXI_GP1_AWVALID),
    .S_AXI_GP1_AWREADY(S_AXI_GP1_AWREADY),
    .S_AXI_GP1_WDATA(S_AXI_GP1_WDATA),
    .S_AXI_GP1_WSTRB(S_AXI_GP1_WSTRB),
    .S_AXI_GP1_WVALID(S_AXI_GP1_WVALID),
    .S_AXI_GP1_WREADY(S_AXI_GP1_WREADY),
    .S_AXI_GP1_BRESP(S_AXI_GP1_BRESP),
    .S_AXI_GP1_BVALID(S_AXI_GP1_BVALID),
    .S_AXI_GP1_BREADY(S_AXI_GP1_BREADY),
    .S_AXI_GP1_ARID(S_AXI_GP1_ARID),
    .S_AXI_GP1_ARADDR(S_AXI_GP1_ARADDR),
    .S_AXI_GP1_ARPROT(S_AXI_GP1_ARPROT),
    .S_AXI_GP1_ARVALID(S_AXI_GP1_ARVALID),
    .S_AXI_GP1_ARREADY(S_AXI_GP1_ARREADY),
    .S_AXI_GP1_RDATA(S_AXI_GP1_RDATA),
    .S_AXI_GP1_RRESP(S_AXI_GP1_RRESP),
    .S_AXI_GP1_RVALID(S_AXI_GP1_RVALID),
    .S_AXI_GP1_RREADY(S_AXI_GP1_RREADY),
    .S_AXI_GP1_AWLEN(S_AXI_GP1_AWLEN),
    .S_AXI_GP1_RLAST(S_AXI_GP1_RLAST),
    .S_AXI_GP1_ARCACHE(S_AXI_GP1_ARCACHE),
    .S_AXI_GP1_AWSIZE(S_AXI_GP1_AWSIZE),
    .S_AXI_GP1_AWBURST(S_AXI_GP1_AWBURST),
    .S_AXI_GP1_AWCACHE(S_AXI_GP1_AWCACHE),
    .S_AXI_GP1_WLAST(S_AXI_GP1_WLAST),
    .S_AXI_GP1_ARLEN(S_AXI_GP1_ARLEN),
    .S_AXI_GP1_ARBURST(S_AXI_GP1_ARBURST),
    .S_AXI_GP1_ARSIZE(S_AXI_GP1_ARSIZE),

    // Misc Interrupts, GPIO, clk
    .IRQ_F2P(IRQ_F2P),

    .GPIO_I(ps_gpio_in),
    .GPIO_O(ps_gpio_out),
    .GPIO_T(ps_gpio_tri),

    .FCLK_CLK0(clk100),
    .FCLK_RESET0(FCLK_RESET0),
    .FCLK_CLK1(clk40),
    // .FCLK_RESET1(FCLK_RESET1),
    .FCLK_CLK2(meas_clk_ref),
    // .FCLK_RESET2(FCLK_RESET2),
    .FCLK_CLK3(bus_clk),
    // .FCLK_RESET3(FCLK_RESET3),

    // Outward connections to the pins
    .MIO(MIO),
    .DDR_CAS_n(DDR_CAS_n),
    .DDR_CKE(DDR_CKE),
    .DDR_Clk_n(DDR_Clk_n),
    .DDR_Clk(DDR_Clk),
    .DDR_CS_n(DDR_CS_n),
    .DDR_DRSTB(DDR_DRSTB),
    .DDR_ODT(DDR_ODT),
    .DDR_RAS_n(DDR_RAS_n),
    .DDR_WEB(DDR_WEB),
    .DDR_BankAddr(DDR_BankAddr),
    .DDR_Addr(DDR_Addr),
    .DDR_VRN(DDR_VRN),
    .DDR_VRP(DDR_VRP),
    .DDR_DM(DDR_DM),
    .DDR_DQ(DDR_DQ),
    .DDR_DQS_n(DDR_DQS_n),
    .DDR_DQS(DDR_DQS),
    .PS_SRSTB(PS_SRSTB),
    .PS_CLK(PS_CLK),
    .PS_PORB(PS_PORB)
  );

   ///////////////////////////////////////////////////////////////////////////////////
   //
   // Xilinx DDR3 Controller and PHY.
   //
   ///////////////////////////////////////////////////////////////////////////////////


   wire        ddr3_axi_clk;           // 1/4 DDR external clock rate (250MHz)
   wire        ddr3_axi_clk_x2;        // 1/4 DDR external clock rate (250MHz)
   wire        ddr3_axi_rst;           // Synchronized to ddr_sys_clk
   wire        ddr3_running;           // DRAM calibration complete.

   // Slave Interface Write Address Ports
   wire        s_axi_awid;
   wire [31:0] s_axi_awaddr;
   wire [7:0]  s_axi_awlen;
   wire [2:0]  s_axi_awsize;
   wire [1:0]  s_axi_awburst;
   wire [0:0]  s_axi_awlock;
   wire [3:0]  s_axi_awcache;
   wire [2:0]  s_axi_awprot;
   wire [3:0]  s_axi_awqos;
   wire        s_axi_awvalid;
   wire        s_axi_awready;
   // Slave Interface Write Data Ports
   wire [255:0] s_axi_wdata;
   wire [31:0]  s_axi_wstrb;
   wire     s_axi_wlast;
   wire     s_axi_wvalid;
   wire     s_axi_wready;
   // Slave Interface Write Response Ports
   wire     s_axi_bready;
   wire     s_axi_bid;
   wire [1:0]   s_axi_bresp;
   wire     s_axi_bvalid;
   // Slave Interface Read Address Ports
   wire     s_axi_arid;
   wire [31:0]  s_axi_araddr;
   wire [7:0]   s_axi_arlen;
   wire [2:0]   s_axi_arsize;
   wire [1:0]   s_axi_arburst;
   wire [0:0]   s_axi_arlock;
   wire [3:0]   s_axi_arcache;
   wire [2:0]   s_axi_arprot;
   wire [3:0]   s_axi_arqos;
   wire     s_axi_arvalid;
   wire     s_axi_arready;
   // Slave Interface Read Data Ports
   wire     s_axi_rready;
   wire     s_axi_rid;
   wire [255:0] s_axi_rdata;
   wire [1:0]   s_axi_rresp;
   wire     s_axi_rlast;
   wire     s_axi_rvalid;

   reg      ddr3_axi_rst_reg_n;

   // Copied this reset circuit from example design.
   always @(posedge ddr3_axi_clk)
     ddr3_axi_rst_reg_n <= ~ddr3_axi_rst;


   // Instantiate the DDR3 MIG core
   //
   // The top-level IP block has no parameters defined for some reason.
   // Most of configurable parameters are hard-coded in the mig so get
   // some additional knobs we pull those out into verilog headers.
   //
   // Synthesis params:  ip/ddr3_32bit/ddr3_32bit_mig_parameters.vh
   // Simulation params: ip/ddr3_32bit/ddr3_32bit_mig_sim_parameters.vh

   ddr3_32bit u_ddr3_32bit (
      // Memory interface ports
      .ddr3_addr                      (ddr3_addr),
      .ddr3_ba                        (ddr3_ba),
      .ddr3_cas_n                     (ddr3_cas_n),
      .ddr3_ck_n                      (ddr3_ck_n),
      .ddr3_ck_p                      (ddr3_ck_p),
      .ddr3_cke                       (ddr3_cke),
      .ddr3_ras_n                     (ddr3_ras_n),
      .ddr3_reset_n                   (ddr3_reset_n),
      .ddr3_we_n                      (ddr3_we_n),
      .ddr3_dq                        (ddr3_dq),
      .ddr3_dqs_n                     (ddr3_dqs_n),
      .ddr3_dqs_p                     (ddr3_dqs_p),
      .init_calib_complete            (ddr3_running),

      .ddr3_cs_n                      (ddr3_cs_n),
      .ddr3_dm                        (ddr3_dm),
      .ddr3_odt                       (ddr3_odt),
      // Application interface ports
      .ui_clk                         (ddr3_axi_clk),  // 200Hz clock out
      .ui_clk_x2                      (ddr3_axi_clk_x2), //300 MHz, not actually x2 for n310 design because of timing.
      .ui_clk_sync_rst                (ddr3_axi_rst),  // Active high Reset signal synchronised to 200 MHz.
      .aresetn                        (ddr3_axi_rst_reg_n),
      .app_sr_req                     (1'b0),
      .app_sr_active                  (app_sr_active),
      .app_ref_req                    (1'b0),
      .app_ref_ack                    (app_ref_ack),
      .app_zq_req                     (1'b0),
      .app_zq_ack                     (app_zq_ack),
      // Slave Interface Write Address Ports
      .s_axi_awid                     (s_axi_awid),
      .s_axi_awaddr                   (s_axi_awaddr),
      .s_axi_awlen                    (s_axi_awlen),
      .s_axi_awsize                   (s_axi_awsize),
      .s_axi_awburst                  (s_axi_awburst),
      .s_axi_awlock                   (s_axi_awlock),
      .s_axi_awcache                  (s_axi_awcache),
      .s_axi_awprot                   (s_axi_awprot),
      .s_axi_awqos                    (s_axi_awqos),
      .s_axi_awvalid                  (s_axi_awvalid),
      .s_axi_awready                  (s_axi_awready),
      // Slave Interface Write Data Ports
      .s_axi_wdata                    (s_axi_wdata),
      .s_axi_wstrb                    (s_axi_wstrb),
      .s_axi_wlast                    (s_axi_wlast),
      .s_axi_wvalid                   (s_axi_wvalid),
      .s_axi_wready                   (s_axi_wready),
      // Slave Interface Write Response Ports
      .s_axi_bid                      (s_axi_bid),
      .s_axi_bresp                    (s_axi_bresp),
      .s_axi_bvalid                   (s_axi_bvalid),
      .s_axi_bready                   (s_axi_bready),
      // Slave Interface Read Address Ports
      .s_axi_arid                     (s_axi_arid),
      .s_axi_araddr                   (s_axi_araddr),
      .s_axi_arlen                    (s_axi_arlen),
      .s_axi_arsize                   (s_axi_arsize),
      .s_axi_arburst                  (s_axi_arburst),
      .s_axi_arlock                   (s_axi_arlock),
      .s_axi_arcache                  (s_axi_arcache),
      .s_axi_arprot                   (s_axi_arprot),
      .s_axi_arqos                    (s_axi_arqos),
      .s_axi_arvalid                  (s_axi_arvalid),
      .s_axi_arready                  (s_axi_arready),
      // Slave Interface Read Data Ports
      .s_axi_rid                      (s_axi_rid),
      .s_axi_rdata                    (s_axi_rdata),
      .s_axi_rresp                    (s_axi_rresp),
      .s_axi_rlast                    (s_axi_rlast),
      .s_axi_rvalid                   (s_axi_rvalid),
      .s_axi_rready                   (s_axi_rready),
      // System Clock Ports
      .sys_clk_p                       (sys_clk_p),
      .sys_clk_n                       (sys_clk_n),
      .clk_ref_i                       (bus_clk),

      .sys_rst                        (~global_rst) // IJB. Poorly named active low. Should change RST_ACT_LOW.
   );


  ///////////////////////////////////////////////////////
  //
  // DB PS SPI Connections
  //
  ///////////////////////////////////////////////////////

  // DB A SPI Connections
  wire cpld_a_cs_n;
  wire cpld_pl_a_cs_n;
  wire lmk_a_cs_n;
  wire dac_a_cs_n;
  wire myk_a_cs_n;

  // Split out the SCLK and MOSI data to Mykonos and the CPLD.
  assign DBA_CPLD_PS_SPI_SCLK = spi0_sclk;
  assign DBA_CPLD_PS_SPI_SDI  = spi0_mosi;

  //vhook_warn PL SPI connected to the PS right now!
  assign DBA_CPLD_PL_SPI_SCLK = spi0_sclk;
  assign DBA_CPLD_PL_SPI_SDI  = spi0_mosi;

  assign DBA_MYK_SPI_SCLK     = spi0_sclk;
  assign DBA_MYK_SPI_SDIO     = spi0_mosi;

  // Assign individual chip selects from PS SPI MASTER 0.
  assign cpld_a_cs_n = spi0_ss0;
  assign lmk_a_cs_n  = spi0_ss1;
  assign dac_a_cs_n  = ps_gpio_out[8]; // DAC select driven through GPIO.
  assign myk_a_cs_n  = spi0_ss2;

  // Returned data mux from the SPI interfaces.
  assign spi0_miso = ~myk_a_cs_n      ? DBA_MYK_SPI_SDO  : // From Mykonos
                     DBA_CPLD_PS_SPI_SDO;

  // For the PS SPI connection to the CPLD, we use the LE and ADDR lines as individual
  // chip selects for the CPLD endpoint as well as the LMK and DAC endpoints.
  // LE      = CPLD
  // ADDR[0] = LMK
  // ADDR[1] = DAC
  assign DBA_CPLD_PS_SPI_LE       = cpld_a_cs_n;
  assign DBA_CPLD_PL_SPI_LE       = cpld_pl_a_cs_n;
  assign DBA_CPLD_PS_SPI_ADDR[0]  = lmk_a_cs_n;
  assign DBA_CPLD_PS_SPI_ADDR[1]  = dac_a_cs_n;
  assign DBA_MYK_SPI_CS_n         = myk_a_cs_n;


  // Default the other control signals (just for now).
  assign DBA_CH1_TX_DSA_DATA = 6'b0;
  assign DBA_CH1_RX_DSA_DATA = 6'b0;
  assign DBA_CH2_TX_DSA_DATA = 6'b0;
  assign DBA_CH2_RX_DSA_DATA = 6'b0;

  assign DBA_ATR_RX_1 = 1'b1;
  assign DBA_ATR_RX_2 = 1'b1;
  assign DBA_ATR_TX_1 = 1'b1;
  assign DBA_ATR_TX_2 = 1'b1;

  assign DBA_MYK_GPIO_0  = 1'b0;
  assign DBA_MYK_GPIO_1  = 1'b0;
  assign DBA_MYK_GPIO_3  = 1'b0;
  assign DBA_MYK_GPIO_4  = 1'b0;
  assign DBA_MYK_GPIO_12 = 1'b0;
  assign DBA_MYK_GPIO_13 = 1'b0;
  assign DBA_MYK_GPIO_14 = 1'b0;
  assign DBA_MYK_GPIO_15 = 1'b0;



  // DB B SPI Connections
  wire cpld_b_cs_n;
  wire cpld_pl_b_cs_n;
  wire lmk_b_cs_n;
  wire dac_b_cs_n;
  wire myk_b_cs_n;

  // Split out the SCLK and MOSI data to Mykonos and the CPLD.
  assign DBB_CPLD_PS_SPI_SCLK = spi1_sclk;
  assign DBB_CPLD_PS_SPI_SDI  = spi1_mosi;

  assign DBB_MYK_SPI_SCLK     = spi1_sclk;
  assign DBB_MYK_SPI_SDIO     = spi1_mosi;

  // Assign individual chip selects from PS SPI MASTER 1.
  assign cpld_b_cs_n = spi1_ss0;
  assign lmk_b_cs_n  = spi1_ss1;
  assign dac_b_cs_n  = ps_gpio_out[9]; // DAC select driven through GPIO.
  assign myk_b_cs_n  = spi1_ss2;

  // Returned data mux from the SPI interfaces.
  assign spi1_miso = ~myk_b_cs_n      ? DBB_MYK_SPI_SDO  : // From Mykonos
                     DBB_CPLD_PS_SPI_SDO;

  // For the PS SPI connection to the CPLD, we use the LE and ADDR lines as individual
  // chip selects for the CPLD endpoint as well as the LMK and DAC endpoints.
  // LE      = CPLD
  // ADDR[0] = LMK
  // ADDR[1] = DAC
  assign DBB_CPLD_PS_SPI_LE       = cpld_b_cs_n;
  assign DBB_CPLD_PL_SPI_LE       = cpld_pl_b_cs_n;
  assign DBB_CPLD_PS_SPI_ADDR[0]  = lmk_b_cs_n;
  assign DBB_CPLD_PS_SPI_ADDR[1]  = dac_b_cs_n;
  assign DBB_MYK_SPI_CS_n         = myk_b_cs_n;


  // For now, default the DSAs to something low-power... is this right?
  assign DBB_CH1_TX_DSA_DATA = 6'b0;
  assign DBB_CH1_RX_DSA_DATA = 6'b0;
  assign DBB_CH2_TX_DSA_DATA = 6'b0;
  assign DBB_CH2_RX_DSA_DATA = 6'b0;

  assign DBB_ATR_RX_1 = 1'b1;
  assign DBB_ATR_RX_2 = 1'b1;
  assign DBB_ATR_TX_1 = 1'b1;
  assign DBB_ATR_TX_2 = 1'b1;

  assign DBB_MYK_GPIO_0  = 1'b0;
  assign DBB_MYK_GPIO_1  = 1'b0;
  assign DBB_MYK_GPIO_3  = 1'b0;
  assign DBB_MYK_GPIO_4  = 1'b0;
  assign DBB_MYK_GPIO_12 = 1'b0;
  assign DBB_MYK_GPIO_13 = 1'b0;
  assign DBB_MYK_GPIO_14 = 1'b0;
  assign DBB_MYK_GPIO_15 = 1'b0;




  ///////////////////////////////////////////////////////
  //
  // N310 CORE
  //
  ///////////////////////////////////////////////////////

  wire  [31:0]     rx0;
  wire  [31:0]     rx1;
  wire  [31:0]     rx2;
  wire  [31:0]     rx3;
  wire  [31:0]     tx0;
  wire  [31:0]     tx1;
  wire  [31:0]     tx2;
  wire  [31:0]     tx3;
  wire  [3:0]      rx_stb;
  wire  [3:0]      tx_stb;
  wire pps_radioclk1x;

  n310_core #(.REG_AWIDTH(14), .BUS_CLK_RATE(BUS_CLK_RATE)) n310_core
  (
    //Clocks and resets
    .radio_clk(radio_clk),
    .radio_rst(radio_rst),
    .bus_clk(bus_clk),
    .bus_rst(bus_rst),

    // Clocking and PPS Controls/Inidcators
    .pps(pps_radioclk1x),
    .pps_select(pps_select),
    .pps_out_enb(pps_out_enb),
    .ref_clk_reset(),
    .meas_clk_reset(meas_clk_reset),
    .ref_clk_locked(1'b1),
    .meas_clk_locked(meas_clk_locked),

    .s_axi_aclk(clk40),
    .s_axi_aresetn(FCLK_RESET0N),
    // AXI4-Lite: Write address port (domain: s_axi_aclk)
    .s_axi_awaddr(M_AXI_GP0_AWADDR_S4),
    .s_axi_awvalid(M_AXI_GP0_AWVALID_S4),
    .s_axi_awready(M_AXI_GP0_AWREADY_S4),
    // AXI4-Lite: Write data port (domain: s_axi_aclk)
    .s_axi_wdata(M_AXI_GP0_WDATA_S4),
    .s_axi_wstrb(M_AXI_GP0_WSTRB_S4),
    .s_axi_wvalid(M_AXI_GP0_WVALID_S4),
    .s_axi_wready(M_AXI_GP0_WREADY_S4),
    // AXI4-Lite: Write response port (domain: s_axi_aclk)
    .s_axi_bresp(M_AXI_GP0_BRESP_S4),
    .s_axi_bvalid(M_AXI_GP0_BVALID_S4),
    .s_axi_bready(M_AXI_GP0_BREADY_S4),
    // AXI4-Lite: Read address port (domain: s_axi_aclk)
    .s_axi_araddr(M_AXI_GP0_ARADDR_S4),
    .s_axi_arvalid(M_AXI_GP0_ARVALID_S4),
    .s_axi_arready(M_AXI_GP0_ARREADY_S4),
    // AXI4-Lite: Read data port (domain: s_axi_aclk)
    .s_axi_rdata(M_AXI_GP0_RDATA_S4),
    .s_axi_rresp(M_AXI_GP0_RRESP_S4),
    .s_axi_rvalid(M_AXI_GP0_RVALID_S4),
    .s_axi_rready(M_AXI_GP0_RREADY_S4),

    // JESD204
    .rx0(rx0),
    .tx0(tx0),
    .rx1(rx1),
    .tx1(tx1),
    .rx2(rx2),
    .tx2(tx2),
    .rx3(rx3),
    .tx3(tx3),
    .rx_stb(rx_stb),
    .tx_stb(tx_stb),

    //DMA
    .dmao_tdata(),
    .dmao_tlast(),
    .dmao_tvalid(),
    .dmao_tready(),

    .dmai_tdata(),
    .dmai_tlast(),
    .dmai_tvalid(),
    .dmai_tready(),

    // DRAM signals.
    .ddr3_axi_clk              (ddr3_axi_clk),
    .ddr3_axi_clk_x2           (ddr3_axi_clk_x2),
    .ddr3_axi_rst              (ddr3_axi_rst),
    .ddr3_running              (ddr3_running),
    // Slave Interface Write Address Ports
    .ddr3_axi_awid             (s_axi_awid),
    .ddr3_axi_awaddr           (s_axi_awaddr),
    .ddr3_axi_awlen            (s_axi_awlen),
    .ddr3_axi_awsize           (s_axi_awsize),
    .ddr3_axi_awburst          (s_axi_awburst),
    .ddr3_axi_awlock           (s_axi_awlock),
    .ddr3_axi_awcache          (s_axi_awcache),
    .ddr3_axi_awprot           (s_axi_awprot),
    .ddr3_axi_awqos            (s_axi_awqos),
    .ddr3_axi_awvalid          (s_axi_awvalid),
    .ddr3_axi_awready          (s_axi_awready),
    // Slave Interface Write Data Ports
    .ddr3_axi_wdata            (s_axi_wdata),
    .ddr3_axi_wstrb            (s_axi_wstrb),
    .ddr3_axi_wlast            (s_axi_wlast),
    .ddr3_axi_wvalid           (s_axi_wvalid),
    .ddr3_axi_wready           (s_axi_wready),
    // Slave Interface Write Response Ports
    .ddr3_axi_bid              (s_axi_bid),
    .ddr3_axi_bresp            (s_axi_bresp),
    .ddr3_axi_bvalid           (s_axi_bvalid),
    .ddr3_axi_bready           (s_axi_bready),
    // Slave Interface Read Address Ports
    .ddr3_axi_arid             (s_axi_arid),
    .ddr3_axi_araddr           (s_axi_araddr),
    .ddr3_axi_arlen            (s_axi_arlen),
    .ddr3_axi_arsize           (s_axi_arsize),
    .ddr3_axi_arburst          (s_axi_arburst),
    .ddr3_axi_arlock           (s_axi_arlock),
    .ddr3_axi_arcache          (s_axi_arcache),
    .ddr3_axi_arprot           (s_axi_arprot),
    .ddr3_axi_arqos            (s_axi_arqos),
    .ddr3_axi_arvalid          (s_axi_arvalid),
    .ddr3_axi_arready          (s_axi_arready),
    // Slave Interface Read Data Ports
    .ddr3_axi_rid              (s_axi_rid),
    .ddr3_axi_rdata            (s_axi_rdata),
    .ddr3_axi_rresp            (s_axi_rresp),
    .ddr3_axi_rlast            (s_axi_rlast),
    .ddr3_axi_rvalid           (s_axi_rvalid),
    .ddr3_axi_rready           (s_axi_rready),


    // VITA to Ethernet
    .v2e0_tdata(v2e0_tdata),
    .v2e0_tvalid(v2e0_tvalid),
    .v2e0_tlast(v2e0_tlast),
    .v2e0_tready(v2e0_tready),

    .v2e1_tdata(v2e1_tdata),
    .v2e1_tlast(v2e1_tlast),
    .v2e1_tvalid(v2e1_tvalid),
    .v2e1_tready(v2e1_tready),

    // Ethernet to VITA
    .e2v0_tdata(e2v0_tdata),
    .e2v0_tlast(e2v0_tlast),
    .e2v0_tvalid(e2v0_tvalid),
    .e2v0_tready(e2v0_tready),

    .e2v1_tdata(e2v1_tdata),
    .e2v1_tlast(e2v1_tlast),
    .e2v1_tvalid(e2v1_tvalid),
    .e2v1_tready(e2v1_tready)
  );

  // //////////////////////////////////////////////////////////////////////
  //
  // Daughterboard Cores
  //
  // //////////////////////////////////////////////////////////////////////

  //vhook_sigstart
  wire aAdcSyncUnusedA;
  wire aAdcSyncUnusedB;
  wire aDacSyncUnusedA;
  wire aDacSyncUnusedB;
  wire aLmkSyncUnusedB;
  wire [49:0] bRegPortInFlatA;
  wire [49:0] bRegPortInFlatB;
  wire [33:0] bRegPortOutFlatA;
  wire [33:0] bRegPortOutFlatB;
  wire rRSP_a_unused;
  wire rRSP_b_unused;
  wire rx_a_valid;
  wire rx_b_valid;
  wire sPpsUnusedB;
  wire sRTC_a_unused;
  wire sRTC_b_unused;
  wire tx_a_rfi;
  wire tx_b_rfi;
  //vhook_sigend

  wire          reg_portA_rd;
  wire          reg_portA_wr;
  wire [14-1:0] reg_portA_addr;
  wire [32-1:0] reg_portA_wr_data;
  wire [32-1:0] reg_portA_rd_data;
  wire          reg_portA_ready;
  wire          validA_unused;

  assign bRegPortInFlatA = {2'b0, reg_portA_addr, reg_portA_wr_data, reg_portA_rd, reg_portA_wr};
  assign {reg_portA_rd_data, validA_unused, reg_portA_ready} = bRegPortOutFlatA;

  //vhook   DbCore dba_core
  //vhook_c aReset ~FCLK_RESET0N
  //vhook_a bReset 1'b0
  //vhook_a BusClk clk40
  //vhook_a Clk40  clk40
  //vhook_a MeasClk  meas_clk
  //vhook_a FpgaClk_p DBA_FPGA_CLK_p
  //vhook_a FpgaClk_n DBA_FPGA_CLK_n
  //vhook_a SampleClk1xOut  radio_clk
  //vhook_a SampleClk1x     radio_clk
  //vhook_a SampleClk2xOut  radio_clk_2x
  //vhook_a SampleClk2x     radio_clk_2x
  //vhook_a bRegPortInFlat  bRegPortInFlatA
  //vhook_a bRegPortOutFlat bRegPortOutFlatA
  //vhook_a kSlotId  1'b0
  //vhook_a sSysRefFpgaLvds_p DBA_FPGA_SYSREF_p
  //vhook_a sSysRefFpgaLvds_n DBA_FPGA_SYSREF_n
  //vhook_a aLmkSync DBA_CPLD_PL_SPI_ADDR[2]
  //vhook_a JesdRefClk_p USRPIO_A_MGTCLK_P
  //vhook_a JesdRefClk_n USRPIO_A_MGTCLK_N
  //vhook_a aAdcRx_p   USRPIO_A_RX_P
  //vhook_a aAdcRx_n   USRPIO_A_RX_N
  //vhook_a aSyncAdcOut_n  DBA_MYK_SYNC_IN_n
  //vhook_a aDacTx_p   USRPIO_A_TX_P
  //vhook_a aDacTx_n   USRPIO_A_TX_N
  //vhook_a aSyncDacIn_n   DBA_MYK_SYNC_OUT_n
  //vhook_a aAdcSync aAdcSyncUnusedA
  //vhook_a aDacSync aDacSyncUnusedA
  //vhook_a sAdcDataValid     rx_a_valid
  //vhook_a sAdcDataSamples0I rx0[31:16]
  //vhook_a sAdcDataSamples0Q rx0[15:0]
  //vhook_a sAdcDataSamples1I rx1[31:16]
  //vhook_a sAdcDataSamples1Q rx1[15:0]
  //vhook_a sDacReadyForInput tx_a_rfi
  //vhook_a sDacDataSamples0I tx0[31:16]
  //vhook_a sDacDataSamples0Q tx0[15:0]
  //vhook_a sDacDataSamples1I tx1[31:16]
  //vhook_a sDacDataSamples1Q tx1[15:0]
  //vhook_a RefClk    ref_clk
  //vhook_a rPpsPulse pps_refclk
  //vhook_a rGatedPulseToPin aUnusedPinForTdcA0
  //vhook_a sGatedPulseToPin aUnusedPinForTdcA1
  //vhook_a sPps      pps_radioclk1x
  //vhook_a sRTC sRTC_a_unused
  //vhook_a rRSP rRSP_a_unused
  DbCore
    dba_core (
      .aReset(~FCLK_RESET0N),                  //in  std_logic
      .bReset(1'b0),                           //in  std_logic
      .BusClk(clk40),                          //in  std_logic
      .Clk40(clk40),                           //in  std_logic
      .MeasClk(meas_clk),                      //in  std_logic
      .FpgaClk_p(DBA_FPGA_CLK_p),              //in  std_logic
      .FpgaClk_n(DBA_FPGA_CLK_n),              //in  std_logic
      .SampleClk1xOut(radio_clk),              //out std_logic
      .SampleClk1x(radio_clk),                 //in  std_logic
      .SampleClk2xOut(radio_clk_2x),           //out std_logic
      .SampleClk2x(radio_clk_2x),              //in  std_logic
      .bRegPortInFlat(bRegPortInFlatA),        //in  std_logic_vector(49:0)
      .bRegPortOutFlat(bRegPortOutFlatA),      //out std_logic_vector(33:0)
      .kSlotId(1'b0),                          //in  std_logic
      .sSysRefFpgaLvds_p(DBA_FPGA_SYSREF_p),   //in  std_logic
      .sSysRefFpgaLvds_n(DBA_FPGA_SYSREF_n),   //in  std_logic
      .aLmkSync(DBA_CPLD_PL_SPI_ADDR[2]),      //out std_logic
      .JesdRefClk_p(USRPIO_A_MGTCLK_P),        //in  std_logic
      .JesdRefClk_n(USRPIO_A_MGTCLK_N),        //in  std_logic
      .aAdcRx_p(USRPIO_A_RX_P),                //in  std_logic_vector(3:0)
      .aAdcRx_n(USRPIO_A_RX_N),                //in  std_logic_vector(3:0)
      .aSyncAdcOut_n(DBA_MYK_SYNC_IN_n),       //out std_logic
      .aDacTx_p(USRPIO_A_TX_P),                //out std_logic_vector(3:0)
      .aDacTx_n(USRPIO_A_TX_N),                //out std_logic_vector(3:0)
      .aSyncDacIn_n(DBA_MYK_SYNC_OUT_n),       //in  std_logic
      .aAdcSync(aAdcSyncUnusedA),              //out std_logic
      .aDacSync(aDacSyncUnusedA),              //out std_logic
      .sAdcDataValid(rx_a_valid),              //out std_logic
      .sAdcDataSamples0I(rx0[31:16]),          //out std_logic_vector(15:0)
      .sAdcDataSamples0Q(rx0[15:0]),           //out std_logic_vector(15:0)
      .sAdcDataSamples1I(rx1[31:16]),          //out std_logic_vector(15:0)
      .sAdcDataSamples1Q(rx1[15:0]),           //out std_logic_vector(15:0)
      .sDacReadyForInput(tx_a_rfi),            //out std_logic
      .sDacDataSamples0I(tx0[31:16]),          //in  std_logic_vector(15:0)
      .sDacDataSamples0Q(tx0[15:0]),           //in  std_logic_vector(15:0)
      .sDacDataSamples1I(tx1[31:16]),          //in  std_logic_vector(15:0)
      .sDacDataSamples1Q(tx1[15:0]),           //in  std_logic_vector(15:0)
      .RefClk(ref_clk),                        //in  std_logic
      .rPpsPulse(pps_refclk),                  //in  std_logic
      .rGatedPulseToPin(aUnusedPinForTdcA0),   //inout std_logic
      .sGatedPulseToPin(aUnusedPinForTdcA1),   //inout std_logic
      .rRSP(rRSP_a_unused),                    //out std_logic
      .sRTC(sRTC_a_unused),                    //out std_logic
      .sPps(pps_radioclk1x));                  //out std_logic

  assign rx_stb[0] = rx_a_valid;
  assign rx_stb[1] = rx_a_valid;
  assign tx_stb[0] = tx_a_rfi;
  assign tx_stb[1] = tx_a_rfi;

  axil_to_ni_regport #(
    .RP_DWIDTH   (32),
    .RP_AWIDTH   (14),
    .TIMEOUT     (512)
  ) ni_regportA_inst (
    // Clock and reset
    .s_axi_aclk    (clk40),
    .s_axi_areset  (~FCLK_RESET0N),
    // AXI4-Lite: Write address port (domain: s_axi_aclk)
    .s_axi_awaddr  (M_AXI_GP0_AWADDR_S5),
    .s_axi_awvalid (M_AXI_GP0_AWVALID_S5),
    .s_axi_awready (M_AXI_GP0_AWREADY_S5),
    // AXI4-Lite: Write data port (domain: s_axi_aclk)
    .s_axi_wdata   (M_AXI_GP0_WDATA_S5),
    .s_axi_wstrb   (M_AXI_GP0_WSTRB_S5),
    .s_axi_wvalid  (M_AXI_GP0_WVALID_S5),
    .s_axi_wready  (M_AXI_GP0_WREADY_S5),
    // AXI4-Lite: Write response port (domain: s_axi_aclk)
    .s_axi_bresp   (M_AXI_GP0_BRESP_S5),
    .s_axi_bvalid  (M_AXI_GP0_BVALID_S5),
    .s_axi_bready  (M_AXI_GP0_BREADY_S5),
    // AXI4-Lite: Read address port (domain: s_axi_aclk)
    .s_axi_araddr  (M_AXI_GP0_ARADDR_S5),
    .s_axi_arvalid (M_AXI_GP0_ARVALID_S5),
    .s_axi_arready (M_AXI_GP0_ARREADY_S5),
    // AXI4-Lite: Read data port (domain: s_axi_aclk)
    .s_axi_rdata   (M_AXI_GP0_RDATA_S5),
    .s_axi_rresp   (M_AXI_GP0_RRESP_S5),
    .s_axi_rvalid  (M_AXI_GP0_RVALID_S5),
    .s_axi_rready  (M_AXI_GP0_RREADY_S5),
    // Register port
    .reg_port_in_rd    (reg_portA_rd),
    .reg_port_in_wt    (reg_portA_wr),
    .reg_port_in_addr  (reg_portA_addr),
    .reg_port_in_data  (reg_portA_wr_data),
    .reg_port_out_data (reg_portA_rd_data),
    .reg_port_out_ready(reg_portA_ready)
  );


  // Default to '1' since these are actually CS_n lines to the LOs.
  assign DBA_CPLD_PL_SPI_ADDR[0] = 1'b1;
  assign DBA_CPLD_PL_SPI_ADDR[1] = 1'b1;

  assign DBB_CPLD_PL_SPI_ADDR[0] = 1'b1;
  assign DBB_CPLD_PL_SPI_ADDR[1] = 1'b1;


  wire          reg_portB_rd;
  wire          reg_portB_wr;
  wire [14-1:0] reg_portB_addr;
  wire [32-1:0] reg_portB_wr_data;
  wire [32-1:0] reg_portB_rd_data;
  wire          reg_portB_ready;
  wire          validB_unused;

  assign bRegPortInFlatB = {2'b0, reg_portB_addr, reg_portB_wr_data, reg_portB_rd, reg_portB_wr};
  assign {reg_portB_rd_data, validB_unused, reg_portB_ready} = bRegPortOutFlatB;

  //vhook   DbCore dbb_core
  //vhook_c aReset ~FCLK_RESET0N
  //vhook_a bReset 1'b0
  //vhook_a BusClk clk40
  //vhook_a Clk40  clk40
  //vhook_a MeasClk  meas_clk
  //vhook_a FpgaClk_p DBB_FPGA_CLK_p
  //vhook_a FpgaClk_n DBB_FPGA_CLK_n
  //vhook_a SampleClk1xOut  radio_clkB
  //vhook_a SampleClk1x     radio_clk
  //vhook_a SampleClk2xOut  radio_clk_2xB
  //vhook_a SampleClk2x     radio_clk_2x
  //vhook_a bRegPortInFlat  bRegPortInFlatB
  //vhook_a bRegPortOutFlat bRegPortOutFlatB
  //vhook_a kSlotId  1'b1
  //vhook_a sSysRefFpgaLvds_p DBB_FPGA_SYSREF_p
  //vhook_a sSysRefFpgaLvds_n DBB_FPGA_SYSREF_n
  //vhook_a aLmkSync DBB_CPLD_PL_SPI_ADDR[2]
  //vhook_a JesdRefClk_p USRPIO_B_MGTCLK_P
  //vhook_a JesdRefClk_n USRPIO_B_MGTCLK_N
  //vhook_a aAdcRx_p   USRPIO_B_RX_P
  //vhook_a aAdcRx_n   USRPIO_B_RX_N
  //vhook_a aSyncAdcOut_n  DBB_MYK_SYNC_IN_n
  //vhook_a aDacTx_p   USRPIO_B_TX_P
  //vhook_a aDacTx_n   USRPIO_B_TX_N
  //vhook_a aSyncDacIn_n   DBB_MYK_SYNC_OUT_n
  //vhook_a aAdcSync aAdcSyncUnusedB
  //vhook_a aDacSync aDacSyncUnusedB
  //vhook_a sAdcDataValid     rx_b_valid
  //vhook_a sAdcDataSamples0I rx2[31:16]
  //vhook_a sAdcDataSamples0Q rx2[15:0]
  //vhook_a sAdcDataSamples1I rx3[31:16]
  //vhook_a sAdcDataSamples1Q rx3[15:0]
  //vhook_a sDacReadyForInput tx_b_rfi
  //vhook_a sDacDataSamples0I tx2[31:16]
  //vhook_a sDacDataSamples0Q tx2[15:0]
  //vhook_a sDacDataSamples1I tx3[31:16]
  //vhook_a sDacDataSamples1Q tx3[15:0]
  //vhook_a RefClk    ref_clk
  //vhook_a rPpsPulse pps_refclk
  //vhook_a rGatedPulseToPin aUnusedPinForTdcB0
  //vhook_a sGatedPulseToPin aUnusedPinForTdcB1
  //vhook_a sPps sPpsUnusedB
  //vhook_a sRTC sRTC_b_unused
  //vhook_a rRSP rRSP_b_unused
  DbCore
    dbb_core (
      .aReset(~FCLK_RESET0N),                  //in  std_logic
      .bReset(1'b0),                           //in  std_logic
      .BusClk(clk40),                          //in  std_logic
      .Clk40(clk40),                           //in  std_logic
      .MeasClk(meas_clk),                      //in  std_logic
      .FpgaClk_p(DBB_FPGA_CLK_p),              //in  std_logic
      .FpgaClk_n(DBB_FPGA_CLK_n),              //in  std_logic
      .SampleClk1xOut(radio_clkB),             //out std_logic
      .SampleClk1x(radio_clk),                 //in  std_logic
      .SampleClk2xOut(radio_clk_2xB),          //out std_logic
      .SampleClk2x(radio_clk_2x),              //in  std_logic
      .bRegPortInFlat(bRegPortInFlatB),        //in  std_logic_vector(49:0)
      .bRegPortOutFlat(bRegPortOutFlatB),      //out std_logic_vector(33:0)
      .kSlotId(1'b1),                          //in  std_logic
      .sSysRefFpgaLvds_p(DBB_FPGA_SYSREF_p),   //in  std_logic
      .sSysRefFpgaLvds_n(DBB_FPGA_SYSREF_n),   //in  std_logic
      .aLmkSync(DBB_CPLD_PL_SPI_ADDR[2]),      //out std_logic
      .JesdRefClk_p(USRPIO_B_MGTCLK_P),        //in  std_logic
      .JesdRefClk_n(USRPIO_B_MGTCLK_N),        //in  std_logic
      .aAdcRx_p(USRPIO_B_RX_P),                //in  std_logic_vector(3:0)
      .aAdcRx_n(USRPIO_B_RX_N),                //in  std_logic_vector(3:0)
      .aSyncAdcOut_n(DBB_MYK_SYNC_IN_n),       //out std_logic
      .aDacTx_p(USRPIO_B_TX_P),                //out std_logic_vector(3:0)
      .aDacTx_n(USRPIO_B_TX_N),                //out std_logic_vector(3:0)
      .aSyncDacIn_n(DBB_MYK_SYNC_OUT_n),       //in  std_logic
      .aAdcSync(aAdcSyncUnusedB),              //out std_logic
      .aDacSync(aDacSyncUnusedB),              //out std_logic
      .sAdcDataValid(rx_b_valid),              //out std_logic
      .sAdcDataSamples0I(rx2[31:16]),          //out std_logic_vector(15:0)
      .sAdcDataSamples0Q(rx2[15:0]),           //out std_logic_vector(15:0)
      .sAdcDataSamples1I(rx3[31:16]),          //out std_logic_vector(15:0)
      .sAdcDataSamples1Q(rx3[15:0]),           //out std_logic_vector(15:0)
      .sDacReadyForInput(tx_b_rfi),            //out std_logic
      .sDacDataSamples0I(tx2[31:16]),          //in  std_logic_vector(15:0)
      .sDacDataSamples0Q(tx2[15:0]),           //in  std_logic_vector(15:0)
      .sDacDataSamples1I(tx3[31:16]),          //in  std_logic_vector(15:0)
      .sDacDataSamples1Q(tx3[15:0]),           //in  std_logic_vector(15:0)
      .RefClk(ref_clk),                        //in  std_logic
      .rPpsPulse(pps_refclk),                  //in  std_logic
      .rGatedPulseToPin(aUnusedPinForTdcB0),   //inout std_logic
      .sGatedPulseToPin(aUnusedPinForTdcB1),   //inout std_logic
      .rRSP(rRSP_b_unused),                    //out std_logic
      .sRTC(sRTC_b_unused),                    //out std_logic
      .sPps(sPpsUnusedB));                     //out std_logic

  assign rx_stb[2] = rx_b_valid;
  assign rx_stb[3] = rx_b_valid;
  assign tx_stb[2] = tx_b_rfi;
  assign tx_stb[3] = tx_b_rfi;

  axil_to_ni_regport #(
    .RP_DWIDTH   (32),
    .RP_AWIDTH   (14),
    .TIMEOUT     (512)
  ) ni_regportB_inst (
    // Clock and reset
    .s_axi_aclk    (clk40),
    .s_axi_areset  (~FCLK_RESET0N),
    // AXI4-Lite: Write address port (domain: s_axi_aclk)
    .s_axi_awaddr  (M_AXI_GP0_AWADDR_S6),
    .s_axi_awvalid (M_AXI_GP0_AWVALID_S6),
    .s_axi_awready (M_AXI_GP0_AWREADY_S6),
    // AXI4-Lite: Write data port (domain: s_axi_aclk)
    .s_axi_wdata   (M_AXI_GP0_WDATA_S6),
    .s_axi_wstrb   (M_AXI_GP0_WSTRB_S6),
    .s_axi_wvalid  (M_AXI_GP0_WVALID_S6),
    .s_axi_wready  (M_AXI_GP0_WREADY_S6),
    // AXI4-Lite: Write response port (domain: s_axi_aclk)
    .s_axi_bresp   (M_AXI_GP0_BRESP_S6),
    .s_axi_bvalid  (M_AXI_GP0_BVALID_S6),
    .s_axi_bready  (M_AXI_GP0_BREADY_S6),
    // AXI4-Lite: Read address port (domain: s_axi_aclk)
    .s_axi_araddr  (M_AXI_GP0_ARADDR_S6),
    .s_axi_arvalid (M_AXI_GP0_ARVALID_S6),
    .s_axi_arready (M_AXI_GP0_ARREADY_S6),
    // AXI4-Lite: Read data port (domain: s_axi_aclk)
    .s_axi_rdata   (M_AXI_GP0_RDATA_S6),
    .s_axi_rresp   (M_AXI_GP0_RRESP_S6),
    .s_axi_rvalid  (M_AXI_GP0_RVALID_S6),
    .s_axi_rready  (M_AXI_GP0_RREADY_S6),
    // Register port
    .reg_port_in_rd    (reg_portB_rd),
    .reg_port_in_wt    (reg_portB_wr),
    .reg_port_in_addr  (reg_portB_addr),
    .reg_port_in_data  (reg_portB_wr_data),
    .reg_port_out_data (reg_portB_rd_data),
    .reg_port_out_ready(reg_portB_ready)
  );


  // //////////////////////////////////////////////////////////////////////
  //
  // LEDS
  //
  // //////////////////////////////////////////////////////////////////////

   reg [31:0] counter1;
   always @(posedge bus_clk) begin
     if (FCLK_RESET0)
       counter1 <= 32'd0;
     else
       counter1 <= counter1 + 32'd1;
   end
   reg [31:0] counter2;
   always @(posedge radio_clk) begin
     if (FCLK_RESET0)
       counter2 <= 32'd0;
     else
       counter2 <= counter2 + 32'd1;
   end
   reg [31:0] counter3;
   // always @(posedge gige_refclk) begin
     // if (FCLK_RESET0)
       // counter3 <= 32'd0;
     // else
       // counter3 <= counter3 + 32'd1;
   // end

   assign {SFP_0_LED_B, SFP_1_LED_B} = {sfp0_phy_status[0],sfp1_phy_status[0]};

   assign PANEL_LED_LINK = counter1[26];
   assign PANEL_LED_REF = counter2[26];
   assign PANEL_LED_GPS = counter3[26];

   // Check Clock frequency through PPS_OUT

   // TODO:  Only for DEBUG
   // ODDR #(
      // .DDR_CLK_EDGE("SAME_EDGE"), // "OPPOSITE_EDGE" or "SAME_EDGE"
      // .INIT(1'b0),    // Initial value of Q: 1'b0 or 1'b1
      // .SRTYPE("SYNC") // Set/Reset type: "SYNC" or "ASYNC"
   // ) fclk_inst (
      // .Q(REF_1PPS_OUT),   // 1-bit DDR output
      // .C(gige_refclk),   // 1-bit clock input
      // .CE(1'b1), // 1-bit clock enable input
      // .D1(1'b0), // 1-bit data input (positive edge)
      // .D2(1'b1), // 1-bit data input (negative edge)
      // .R(1'b0),   // 1-bit reset
      // .S(1'b0)    // 1-bit set
   // );

endmodule
