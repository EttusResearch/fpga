
// Copyright 2014 Ettus Research

// Assumes 32-bit elements (like 16cs) carried over AXI
// User block controls packet sizes with tlast
// simple_mode=1 allows user to ignore chdr stuff, must produce 1 packet for each one consume
// simple_mode=0 user controls all chdr info, must control s_axis_data_tuser

// _tuser bit definitions
//   [127:64] == CHDR header
//   [63:0] == timestamp

module axi_wrapper
  #(parameter BASE=128,
    parameter NUM_AXI_CONFIG_BUS=1,
    parameter CONFIG_BUS_FIFO_DEPTH=5,
    parameter SIMPLE_MODE=1)
   (input clk, input reset,

    input clear_tx_seqnum,

    // To NoC Shell
    input set_stb, input [7:0] set_addr, input [31:0] set_data,
    input [63:0] i_tdata, input i_tlast, input i_tvalid, output i_tready,
    output [63:0] o_tdata, output o_tlast, output o_tvalid, input o_tready,
    
    // To AXI IP
    output [31:0] m_axis_data_tdata, output [127:0] m_axis_data_tuser, output m_axis_data_tlast, output m_axis_data_tvalid, input m_axis_data_tready,
    input [31:0] s_axis_data_tdata, input [127:0] s_axis_data_tuser, input s_axis_data_tlast, input s_axis_data_tvalid, output s_axis_data_tready,
    
    // Variable number of AXI configuration busses
    output [NUM_AXI_CONFIG_BUS*32-1:0] m_axis_config_tdata, 
    output [NUM_AXI_CONFIG_BUS-1:0] m_axis_config_tlast, 
    output [NUM_AXI_CONFIG_BUS-1:0] m_axis_config_tvalid, 
    input [NUM_AXI_CONFIG_BUS-1:0] m_axis_config_tready
    );

   // /////////////////////////////////////////////////////////
   // Input side handling, chdr_deframer
   wire [127:0]  m_axis_data_tuser;
   
   chdr_deframer chdr_deframer
     (.clk(clk), .reset(reset), .clear(1'b0),
      .i_tdata(i_tdata), .i_tlast(i_tlast), .i_tvalid(i_tvalid), .i_tready(i_tready),
      .o_tdata(m_axis_data_tdata), .o_tuser(m_axis_data_tuser), .o_tlast(m_axis_data_tlast), .o_tvalid(m_axis_data_tvalid), .o_tready(m_axis_data_tready));

   // /////////////////////////////////////////////////////////
   // Insert time and burst handling here.  A simple FIFO works only if packets are produced 1-for-1 (they may be of different sizes, though)
   wire [15:0] 	 next_destination;
   wire [127:0]  s_axis_data_tuser_int;
   reg 		 sof_in = 1'b1;

   always @(posedge clk)
     if(reset)
       sof_in <= 1'b1;
     else
       if(m_axis_data_tvalid & m_axis_data_tready)
	 sof_in <= ~m_axis_data_tlast;
   
   generate
      if(SIMPLE_MODE)
	begin
	   // Set next destination in chain
	   setting_reg #(.my_addr(BASE), .width(16)) new_destination
	     (.clk(clk), .rst(reset), .strobe(set_stb), .addr(set_addr), .in(set_data),
	      .out(next_destination[15:0]));
	   // FIFO for 
	   axi_fifo_short #(.WIDTH(128)) header_fifo
	     (.clk(clk), .reset(reset), .clear(1'b0),
	      .i_tdata({m_axis_data_tuser[127:96],m_axis_data_tuser[79:64],next_destination,m_axis_data_tuser[63:0]}),
	      .i_tvalid(sof_in&m_axis_data_tvalid&m_axis_data_tready), .i_tready(),
	      .o_tdata(s_axis_data_tuser_int), .o_tvalid(), .o_tready(s_axis_data_tlast&s_axis_data_tvalid&s_axis_data_tready));
	end // if (SIMPLE_MODE)
      else
	assign s_axis_data_tuser_int = s_axis_data_tuser;
   endgenerate
   
   // /////////////////////////////////////////////////////////
   // Output side handling, chdr_framer
   chdr_framer #(.SIZE(10)) chdr_framer
     (.clk(clk), .reset(reset), .clear(clear_tx_seqnum),
      .i_tdata(s_axis_data_tdata), .i_tuser(s_axis_data_tuser_int), .i_tlast(s_axis_data_tlast), .i_tvalid(s_axis_data_tvalid), .i_tready(s_axis_data_tready),
      .o_tdata(o_tdata), .o_tlast(o_tlast), .o_tvalid(o_tvalid), .o_tready(o_tready));

   // /////////////////////////////////////////////////////////
   // Control bus handling
   // FIXME we could put inline control here...
   // Generate additional AXI stream interfaces for configuration. 
   // FIXME need to make sure we don't overrun this if core can backpressure us
   // Write to BASE+8+2*(CONFIG BUS #) asserts tvalid, BASE+8+2*(CONFIG BUS #)+1 asserts tvalid & tlast
   genvar k;
   generate
      for (k = 0; k < NUM_AXI_CONFIG_BUS; k = k + 1) begin
         axi_fifo #(.WIDTH(33), .SIZE(CONFIG_BUS_FIFO_DEPTH)) config_stream
           (.clk(clk), .reset(reset), .clear(1'b0),
            .i_tdata({(set_addr == (BASE+1+2*k+1)),set_data}), .i_tvalid(set_stb & ((set_addr == (BASE+1+2*k))|(set_addr == (BASE+1+2*k+1)))), .i_tready(),
            .o_tdata({m_axis_config_tlast[k],m_axis_config_tdata[32*k+31:32*k]}), .o_tvalid(m_axis_config_tvalid[k]), .o_tready(m_axis_config_tready[k]));
      end
   endgenerate
   
endmodule // axi_wrapper
