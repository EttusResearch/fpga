//
// Copyright 2019 Ettus Research, A National Instruments Company
//
// SPDX-License-Identifier: LGPL-3.0-or-later
//

// Add all new transport types here
localparam [7:0] NODE_TYPE_XPORT_GENERIC = NODE_TYPE_XPORT_BASE + 8'd0;
